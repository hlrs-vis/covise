MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       �:Á�[�҆[�҆[�ҏ#8ү[�ҏ#.�[�ҡ��҅[�҆[���[�ҏ#)��[�ҏ#?҇[�ҏ#<҇[��Rich�[��                PE  L 6ڀL        � !	  �       ��                                                              �8 [   � (                            � �g  `                                            T� ,                          .textbsszl                        �  �.text   I�  �  �                   `.rdata  +*    ,  �             @  @.data   �L   @  $   �             @  �.idata     �     �             @  �.reloc  *y   �  z   �             @  B                                                                                                                                                                                                                                                                                                                        ������ �  �( �H �|
 �  �x� �! �ޛ	 �9� �% ��c �z ��5 �D �[�
 �֧
 ��� �,� ��& �"� ��� �H �% �>� �9� �� �� �*� �� ���	 � �C �!= �\� �G� �� �=� �h�
 �a �� �i� 鴐 �O� ��	 �" ��C �� ��e 顛 �� 釆 �8 �M�
 鸋 �F �� 鉤 �� ��  ��	 �t ��  ��� �� �o �s ��
 �[ �M�
 阄 �c� ��! �/ ��< �� �z� �U� �  �+6 �� �!� �| 采 �"� �J �h� �Ӂ ��X �D �t� �_� � �s �0g �q � �� �<� ���
 �d ��
 ��y 鳅 �nk �i� �� �� �i �� � �+� 香 �q� �<� �� �d �� � �CX �N� �9 �t �) ���  鵩 ��� �k �&7 �A� � ��� ��� �m�	 �� �#<
 �I ���  �4�	 �� �"	 ��	 � 8 �+4 鶃 �A� �<� �1 颖 �~ � �#� �� �� �� �O= �t
 �_ �� �� �6� �� �U �5 �j
 �y �� �� 鮎 �� 鴊 �/� ��� �K �9 鋠 �* ��: 鼖 �w�  �"8 �} �_ 铊 �>�	 �� �Z �o�  �� � �0 �k�  �V� ��� �d ��� �" �Ͱ ��� ��� 鞨 陓 �� ��9 ��Y ��
 �m
 �k 閧 �A�  ��� �W� ��u �-� �	 �S� ��x ��2 �t �� �j� �%h �0f 黭 �} �A� ��  �} �� �] �8� �C� ��� �I� �� �?� �j� �� �`@ �[ �v� ��� ��� ��	 ��g �� �x	 �S@ �n� ��m 餫 �:� �� ��! �P� ��( �V� ��T
 �܇ ��p �1 �M �xC �S� 龽 � �D* �)	 �z� �J �� � �v} �Q3 �|l �4 ��� �=5 �h� �c� �N�  �� �K
 �ߌ
 �j� �� �@� �_
 ��	 ��� ��} �q ��= �-� �y �3� ��
 �1 �@ ��}
 �
6 �� � �K� �F� �q� ��{ �G �rR �� � �� �| ��# �$� ��� ��
 �E~ �З ��� �6d �Q! �� �7� �rC ��7 �8� �C� �NV �i� �TF 鏑 �ڌ
 �E
 �p} �} �� �A� ��� 駅 �� � �� �� �N ��| �2 �� � �u% �@�  �` �V! �AY ��[ �� �� �� �� �Sa �N� �ih
 �t�  �� � �% � ��  �� ��  �j �W� �� �a �H�  �3� �> �y� �$' �� �j �� ��: �n �� �1~ �lc
 �\ �r� �}} �x�  �s� ���  ��� ��v �� �� �U�	 頼 �a �6 �a	 �� 釣 ��I �-�	 � �� �N� �Yg �t� ��w �h � ��� �{O 鶐 �� �g ��	 �Rs �_ �W � �.2 ��: �ԍ �8 ��8 �e� �@? �[W �֖  �!� �' �, ��T ���	 �(�	 ��2 �/ �� �Ԣ �� � � ��n �[� �p �1� ��D �g �t �� �Xn �S �n� �� ��;	 �/  �Zb �%6 �@� � �} �a�
 ��� �7�	 �bD 鍑 �- �" � �: �V �/� �:� ���	 �M � ��� ��C �� �gx
 ��	 �� 鈧 �S ��& �	j	 鴯 �� �� ��� ��� ��g
 ��:	 �12 �= �F ��  �\ �K �c� 鞎
 �g
 �� ��  �  �  �p� �� �F. ���  �  ��` �b; �]/ �, 飁	 ��~ �~�	 餈 �/4 �*� �%�	 �P� �ۧ �" �! �| �ȹ	 � ��] �� �#� ��  鹑
 ��$ �� � ��? �PN ��
 �( �A�	 �lj	 �� �� 魐 ��& �Cy �^�	 �Yv	 ��� �� �� 饝 ��	 �� ��� ��� ��0 �x �2� ��� �h� �' ��T �y= �t� �% �zU �% �0I �8 ��
 ��d
 ��
 � � �Mf �8� �� �^� �) �T  �O� �Z� �B	 �  �s � � �,i �� �R� �� �x� �� �^s �)�  �$� �� �� � ��� ��X �N �Q~ �� �7� ��� ��h �h� 铞 �M 鉤  ��� 鿈 ���
 �f ��  �{� �j �� �,� ��� �B� ��  ��� �s �n� ��� �t' �) �
� �� � J � �' �AU �� �7q �R{ �-� �X� �� �^� �v �t�	 �� �� �! �@� �� �� �A^
 �D ��Y
 �n �G �ع ��A
 �� ��V �H �߂ �*t ��� ���  �4 ��� �qe �U �' �bg 魧 騷 铋 �� �Ix  �$� �Z �ڂ ��� 速 �� �f~ �q{ ��� �w ��	 ��� �� ��V �� �� �T� �/� �� ��� �P: �;D �v) �N
 �� �W� ��} �=�  �8v
 �s� � �ٶ � �/	 �z�  �Eq ��� �k� �M ��	 �� �5 �2� ��" �H� �z �>[ ��� �j �� � �@� �� ��� ��v ��  ��| ��. 颅	 � ��| �, �^� �O ��F ��� �* ��j �� ��
 �f ��� �	 �+
 ��� � �� �v ��  �) ��� �e 骹 �5% ���
 �� �6 �m�
 �,� �� �� �]� 鈎  �3� �� �� ��t
 �?� �z? �e�
 ��* � �� ��" �� �7M �"Y	 �� �x� �Û ���	 �� �T] �_U �:� �_ �P� ���  �� 鱾 �L^ �� �  ��x �H	 �C) � ��  �t� 鏂 �:h �e ��; 黂 馁 �� �/ �� 钄 ��q ��{ ��� �΅ ���	 ��` �O� �< �# �0V �+h �0 �� �� ��� ��0 靖 ��N �v �nK �9� �� �� �H �e� � ) �� �f �ѡ �L� �7* �R�  �� �xM �C�	 �n]
 �� �t� �x  �
� ��> �P� �;# �F� �� ��  �� �"� �� �D �o � ��_
 �� ���
 隙 �u� ��G �� ��< ��K �,� �g� �B� �]� �h �CA 龥 �+ �1 �
 ��- �� �p� ��� �F] �a�  � �'� �� � �s 鳓 �� �)^ �4� �oi �� ��z ��� �� �� �� ��X
 ��� �� ��� �(o
 �c^
 �� �)� �� ��� �B �� ��w �� ��	 �A� �l: �� �2$ � ��� ��j �S ��> �i �?s �*� �Ņ ��n
 �+� ��b �� 鬏 �w� ��� � �8S � �: �Y� �5 �� ��H �5* �  �+C �FW
 �q �� �v �": 鍝 鈮 �s� �p�
 �y� � �o�
 骿 �%� � �6 �� ��! �t �� �& �}� ��  �m �� �y� ��  �� �Z� �%� �^ �K�
 ��c �a �� ��: �2� ��M ��; �n
 ��� ���  ��'
 韩 �:N �� �\ ���  �v9 �; 鬮 ��� �� 魣 ��  �ì  �ޟ  ��Z
 �d 鿅
 銙 �A 骺 �� ��  ��n �� �'�
 �� �=s  �+ 飆 �E �. �Y
 �_� �� �eB ��n
 �kE ��m
 �q� � ��P 鲂 � �a
 �3� 鞺  �l �L�	 ��2 �ڰ �e �@� �� ��	 ��� �<a
 �7� �Җ �ݔ ��0 �30 ��� � �4� � 麉 �� ��U
 �+} �l �� �� �' �2p �T �X4 �#, �� �ij 鴧 �k �
w �U� �`?	 �K� �� �A� �� �g0 ��? �]� ��m � �^! ��
 �To �� ��� ��G �0! � �6� �ѣ �~ �G� ��_ �M� �ؚ �z �~� 鉿 �$� 鏍 �� �� ��� �{u �o �I �L� �G� �S �M� �H� ��{  �~& �)�  ��� �� ��� �� �� ��� ��	 �1� 霶 �7� ��^ �mZ
 ��� �t �� �Iq �4� �?� �z�  �Eu �Pv �2 �&1
 鱆 �� �ט ��� ��� ��  ��� 龯	 �Z ��t ��e ��T
 � �� �+ �6� �х �� ��, �b� 齗 �m �#] � ��� ��~ �� 骷 �e � � �[r �6m  �k 錿 �k �Rg ��- �ع	 � �.� �i> �T0 �L �J�  �U �� ��4 馫 �q�  ��  �� �B_ �t ��� �c� �> ��
 �=	 �ό 骬 �e � � �K� 鶠 ��[
 �� �w0 ��	 �f �z	 �� �Z �)  �D� ��� �
h �En �`z �` �f8 �� �� �U �BZ �{ ��� �#�  �~x  �y �$k �/p �JF �U� ��� 雏
 �&� �A�  �<� �w� ��� �� �� 飑 �� �i� �d� �O� �j� �� � + �- �F �`
 �\O �ǳ �b�	 ��< �� �Ö 鞺 �� 餉 �# �:s �uS �0� �[o �6� �� ��Q �w4 �Rv �A �. �s� �Π	 �)� �� ��I �
y ��� �@v �k� �F[ �AV
 ��> �w �R� � 鸜	 �c ��K �i� ��� �� �J� �%~ ��~ ��� �v�	 �!� 錃 �'E ��/ �}� 阞 �S� �n� �� �z
 �m
 �J� �Š 通 �{7 �5 ��h �|' �׃ ��
 �MO � �c� �>R �I� �Z
 �= �Z �U�  �r �Kg ��� �!\ �<j �G& �p �-* ��	 �M �~. �9&	 �� �3 �jj ��� �p; �� �� �/ �\� �g� ��9 �} �X� �j
 �~� �A �� �ϟ  �� � �@� ���
 �V�	 �1 �\T �'�  �'� �mS �hd �� ��z �y�  � �  ��� �E& �� �b
 馨 �J �<� 駔 ��
 ��`
 �x" �c� ��� ��� � �o	 �� �u� ��? � �v� �;	 ��X �w�
 �x�
 �=� �a ��� �� � �X �6 � ��� ��� �ۉ �� �=	 �|� �w� ��< ��x �� �u �~ ��  餰 ��� �j& �� �� �z ��f �q� �l�  �g�  �p  �� ��� ��  �, �)� �$d ��^	 �Z� �uX �0H �k/ �S �1� �< �� ��x �-� �x� �~	 �� 鹨 ��� �g ��� �" �P �� ���  �!>	 ��
 ��	 ��� ��  �� �c� �� ��� �4� �h
 �:�
 镦	 �$ �+t �� �Q�  � �k
 ��0 魓 騰  ��S
 �� �� ��S �?� �9 �� ��; �` ��. �q 錃 �'�	 ��	 �M� �0 �C�	 ��� �C �� �� ��	 �u� � B ���  �n
 �!� �� �� �r  ��  �� �S� ��� �y� �� �?� �� �eg ��A �[�  �R
 �A ��u
 ��� �B� �m�  ���	 �3	 �3 �I� �dy �_ �� 饁 �p� 雐 ��A �F ��0 �g� �e �={ ��V ��c �� �Y� � �_K ��	 ��i � �;� �V� �!	 � �� �B	 �� 鈱 �$
 �N/ 驸 ��� ��^ 隒 ��� �D 雱	 � �am �̙ �w� �r� �w �� �S� �Ng �F �` �ߋ �[ 饱	 ��. �Y �f� ���  �| �w �b�  �ݞ  ��  �3�
 �n� �: �" ��  �*�	 �p	 �@�	 �} 馄 �a� �v �7t �r� 魰	 ��
 ��� ��� �	q �t
 �^ �Z� �5� �P� �� ��� �> �|m 釸 �d
 ��
 �8| �# �^O �� �m ��  �J � ��� ��q �F�  �1�  �� �W� �m �� �� �S� �  �  ��  ���  �J�  酲 �@� �;b �� �� ��f �wv �r� �=� �( �S�
 �^ �� �t� ��� �J� � �@4	 ��� �z �!p	 霽 �'�  ��� �M� �(�  �6 �d  ��{ �Ā �� �*� ��� ��� �K� �� ��� �|? �g �r �m2 �� �� � 陮 �� �� �[ 镋 �p/ �{�  ��i
 遂 �̳
 ��	 鲭 �= ��� �C �� �I�	 �4	 �k� �[ �� � � �;( �fj  �� �� 闠 �27 ��S �$ �  �.�  � �� ��  �J8 ��
 �0�
 雨	 �vk ��
 �� �7; �", ��
 ��} �s� ��o ��� �Ļ
 �/T ��n �� �pe �� �5
 �1�  ��� �� ��0 ��? �x	 �c_ ��# ��� �( ��  �O �I �P�  ��� �U �� �A �� � �=� 阪 � 鮕 �iC �� �߶ 麔
 �j� � f �� �6�	 �A� �\ 釯 ��  ��� ��E �� �N_ �� 鄁 ��N �j� 饞 �� �;� �V� �1u �n �7f �>	 �r ��8 �� �>� �i�  �Tg �O�  ��� �u ��� �� �V� �ay �<� �W_ �u
 �F
 �>r ��p �ު �y� �Tv �Oc �z{ �et �� �b �� �q �L	 �w9 �b� �-�  ��� �#e �Φ �w  �4` ��a �� �5< � � ��( � ���
 鼦 �� ��T �d  �E �� ��m �	 �� ��� �T� �U� �P�  �+b
 �j� �1� ��F �� �« ��Y �ț �á �^M ��d 鴚 �_A �� �Ō  �6� �k� ��� �� �<� �� ��_ �M�
 �8I �c� �� ��� �� � �j � �`m � �-
 �! �$ �g�  ��o ��; �	 �i �. �	 餺 � ��� �� �p� �Ko �` �� �D �wo ��� �m� �� �S4 ��c �G� �$� �� �Z� � � �  �{^
 ��� �� �� �* �� �m3 �(�
 �d
 �N�  �)n �T� �� �t
 �U9 �@_ �;J �� �� �� �7� ��� �m� �(� �s8 �� �i� �ķ  �X �q
 ��m
 �B �# �C ��� �l� �g� �
 靻 �X �#� �.B �)_ �; �?� �z� �� ��	 �� �f*
 ��+ �l�  � �2/ �I
 �X8 �SX �n�  �l 鴪 �f ��Q ��  �k
 ��_ �vk �!W �|� �w 邽 魿 �| �3�  龊 �9� � ��
 �Z � �`� �o �&L ��  �c	 ��  ��� ��
 �o
 ��	 ��	 �y� �t� �e 銦 ���
 ��m
 �  �ƭ  �a� �Z �{ �r �m{
 ��w �y �p 鉽	 �n �/�  �� �Z �@� �+� �} ��� �� �7�	 �� �=�
 ��� ��C �H
 �L �t�	 �; 隠  配 �@w �C� �F{
 �Q �0� �w �� �s � �� ��  �m
 �% �k 隿	 ��' � �
 �� �k �QJ �|q �ׄ  �[
 ��  �� � �~� �IU �R �o� �Jg ��� � 5 ��X �V�  � ��# �G� �R� ��l
 騿 �#� �� �� ��� �?g ��� ��x � � �� �&l �� �<" 駑 颽 �= ��� ��i �>" �ɒ � ��?
 ��B �- �  鋰 �� �A
 �,! �W �"� �-� 鈿  �C� �4� �9� ��n �P ��k �� � � �{� �G �a� �� ��	 �r� ��� �� �k �� �)� �$� �ϗ �: �� �Е �� �&�	 �, ��H
 �7	 �� �� �: ��  ���  �9i �t� ��	 �	 �E� �`�
 �� �� �< �|\
 闦 �b� ���  �� �Cb ��Q	 �. �t@ �� �� �	 ��h �˒
 �d �ax �<J �7 �R\ �mQ ��� �� �� � �t �/� �0� �j
 �p� ��  �& �W
 �\ ��� �� �m
 �( �3�
 �~�	 �9! ��	 �� �Z� �� �\
 ��I �i ��� ��q
 �W$ �"� ���  ��� �, 鞱 �� �4! 鯡 �*i �Uo �0 �k� �> 遧 �<0 �� �2�  �], �X) �S� �� �yE 鴎 �\ �� � �0 ��r �&q  �4 �^ ���  鲛  �	 �H ��� ��v
 �� �� �� �Z�
 ��	 � �q  �v� �� �� �� ��� �	 鈫 �� ��e �9D �T�  ��� ��� �u�  �@� �0 �� �q@ �l	 �� �� �-� ��s �� ��� �y	 �� �� �:� 饭 ��� �� �� � �^	 �� �� ��m � �3� ��
 �Y� ��� 鿮 骁 ��� �w �KJ �v� �p ��	 �7n ��> ��  �8" �c< �ζ �* �4� �� �� �5Y �Щ 髐 �� ��� �l�  ��� �B
 �� ��g �� ��T ��b �D ��  �
<	 酵 �`) �{$ �@ �A �} �'r �� �m5 �8U ��	 �Μ	 ��) �
 �} ���  鵋 �@x ��\ �v ��j �y �w� 還 �	 �x� �]	 �ީ 鹩 ��~ �_ �jS �%� ���  �+; �ơ  �!P �̒ �� �� �m� ��~ �s1 鮕 �^  �T^  �Y ��? �%A
 �A ��� ��
 ��v ��� �W� �R� ��}
 �n ��: ��� �)�  �$� ��S �:, � �� ��= �V`  �q� �� �p� ��I �m� ��_  �c� �>l �& �Tb �{ �ZQ �U� ��� �& �� �� �|X  ��� � �] 阴 �`  ��5 �Y� 餮  ��� �j| �� ���  雩 �&~ �> �\�	 �ק �L �_
 �, �3� �^� �y) ��U
 �� ��� �u� �`( �+� �� ���
 �z �g� ��* ��� �, �_ � �� ��R ��
 �� �%� �@
 ��5 �m
 �P �l� �7� �B� �� �x� �#�  �� �)Q �dS �1 ��  �g
 ��f �O �[  �Q� �� ��� �� �-	 �� 铳  �c �	� ���
 �o- ��O �5� 鐲
 �[U
 �Vy �� �l ��m  �^� �T �x ��= ��� �Y� �4� �?S ��1 �L ��� �h �&� �A� �L{ ��� �2] ��� 阐 �Ӈ �� �) 鄞	 �N �� �� �p�
 �k� �&� ��� �� �g� � �}� �H� �� �ޠ �� �~ 鯻 �z| �U� �0R �A ��� �1F �Z �׹ ��( ��t � �0 �^> �y, 餠 �% ��w �EY �@� �� �6o ��  �\�  �u �R  �-�  �� �X ��
 驦 �t  鏶 �*�  �]� ��
 �U �2 �A� �<Y ��� �� ��h �9 ��  ��� �	a �+ ��� �N
 � �� ��Q  �� �a� ��` �7� ��P �m� �8� �s �� �i� �| �O� �� �L �� �� ���	 �~ �p� �ǌ ��� �c
 �h� 郘 �� ��\ �t� �x �L �u� �0� �;� �6U �!�  ��6 ��  �� 靎 �(<
 �sT �� �T  �8� �?&	 �ڦ �%� � � ��R �f ��  ��= �WQ ���  �ͣ  �Hd
 �� �α �Y' �Գ �� �ڄ ��  ��	 �' �6� �! ��k �7� �� �8	 �a �S� �.d ��' �t�
 ��	 ��� �� ��� ��� �V� � �̒	 ��� �2�  ��E 鸆 �ñ �h
 �I �4 �T �jK ��	 �l ��N �6 �q� �	 �G� �3 �=�  �he
 ��b	 �V �iM
 �D9 �O� �9 �%� ��� �k� 馦 顃	 �� �'�
 �� �=%	 �� �ӧ �n� ��s 鴸 �� �n� �e� �� ��;
 �F� ��^ ��= �Q �� ��� �ȓ
 ��� � �� ��� �; 骉  �Ş	 ��` ��  �V� �� �܆ ��t �� �� �x �^ ��=
 � �d� �?� �r ��r � a �� �f�  �!� �,� �w� �X �-� �XC �c= �� �Y�
 �� ��  ��Z �
 ��� �; �&R �� � �w� �2B �mF ��� �t �NZ �ٌ	 ��U ��� �*� ��� �P� �6 �6� �� �+ �7�  �. �]& �� �s� ��4 �9 �D� �_� �*( �E�	 ��J � �&� 鑭 ��M �'� ���  �v  �H� �3 鎵  �	H �� 鿰 �� �%� � �� �\ ��; 録
 ��� �� �͘ �Xe  ��� ��� �� ��O �f �� � �0A ��u �&� �� �z �� �� �M� �؇  ��� 龳 �I� �tP �_j ��5 ��� �E �+~ ��y ��m �\� ���  邨 �-� �x� �CN �Α �, �dU �� �
{ �Z 鰤 � �֤ �AN �� �� ��
 ��� �� �q �: ��� �tM 鯂 �: ��* �0� �Z �� �1� ��� �'�	 ��: � �� �C8 �.0 �YP 餆 ��� �y �%g �0� �Z ��K �� �Z �m� �b= �� ��+ ��e
 �� 鹲 �} �O� �� �\ �  �7� 馴 �Av 錴 �7^ �� 靳 ��u ��� �N] �  �T� �_�  �J� �5Y � = �@ �FX �� �,�	 �G� �r} �=� �/ 郏
 鎮  ��5 � �
 �� ��G � � �@ �֞	 ��� �,� �'E ��t �m9 �8K �� ���
 �� �Tb  �O� �Z�	 �� ��� � �&� �r �<�
 ���  �H �}2 �- �#� ��X � �D�  �_� �p ���  ��, � ��l �Ѳ �\� �8
 ��� ��� �, �R �>R
 ��q ��� ��G ��� �5� �P� ��U �`� �� �� ���  �rZ �-� ��� �| �H
 �Y�  ��' ��4 �Z� �U\ � Z ��a �V� �� �Y
 飈	 ��j �< �X8 ��  �>} �6 養 ��� �@ ��G
 �� ��Z �V 遚	 �<� �� 颁 ��' �x� �Ò ��� �� �4� �9 �z� �g �pJ
 �K�	 �` ��� �# �W� �� �-�	 �8? �#C ��} �K �� �� ��; �u= ��G �[W ��	 �� �<� �g? ��� �� ��� �C�
 ��� �� �D �� �ڶ �e�  ��  ��# �6B �� �LZ �WE �2� ��* �tY ��R ��  陞 �$� �o; 骤 �%' �� �K? ��, ��� 霃 ��( �b7 �� �* �S� �.� ��A ��
 ���	 �j�
 ��
 ��� �+2 �Vv ��? �L� ��� �  �]a 鸛 ��& �|	 �� ��Y
 �o� ��n �	 鐩 �+� �F�  �Ѧ
 ��L �G �U �}� ��� �C� �.� �� ��,
 �ߙ	 �~ �Ł � ��� �6� �a�  ��n 駴 �P 靚 �ؔ
 �# ��z ��s �� �o�  �j� �u� �� ��� ��� �m� �L� �� 邎 �mz �� �S�  � �y ��� �o{	 �jz	 酒 � �K �v� �Q� �\4 �� �r�
 �8 �� �� � �� �� �oS �zo �5 � 黵 �6� �q
 �� �g
 �Y
 ��k �HD
 �3� �n� ��	 �$M	 �ϕ �* 镁 鐠 �� �&� ��{ ��
 �j �2F �H �� �� �n4
 �g� ��X	 �Q� �:� �u_  �@� 黋  馃
 ��� �L� ��I �R� ��; �� �� �N9 �ِ �* ��� �� �E� 选 �;� �f�  �Ai �\~ �x	 �2X �=*
 �� ��8 �� �i/ �TZ
 �O �j� �� � B
 �y	 �6  �A� ��� �� �� �&� �hA �� �>! ��P
 �L �� �Z� �U�  �? �~ 鶯 ��r
 �<� ��� �� ��o ��� �#C
 鮵 ��� ��  �G ��n ��� ��b �� �v� �v ��� ��% ��	 ��� 鸣 �sO  �^� �y� �4 �� �Z� �� ��p �+� �f� ��n �O �g� �"� �}� ��� �C	 �� �� �; ��  �:� �� �P� �{P �� ��4 �\� 鷢 �2> �]�	 �(� ��q �� �Y�	 �Z ��Z	 �~ �u ��� �[� �FT �� �	 釳 ��	 �m�	 �q �� �Δ �i� ��� ��  �@� ��& �Л ��@ �� �Q� �\2 �7" ��E ��� �8�
 ��
 �W �i� �t �� ���  ��� �0�  � ��~ �AT �=
 �+ �Bv	 靼 ��� �s� �q ��� � �?w �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������蝺����u3��跢����u3���}�����u3���   _^[���   ;��f�����]�����������������������������������U����   SVW��@����0   ������_^[��]������������U����   SVW��<����1   ������E��<�����<��� t$��<���t� ��c��~����u3���   �	�   �3�_^[���   ;�裑����]��������������������������������U��j�hΡd�    P��8  SVWQ�������N   ������Y�XD3ŉE�P�E�d�    �M�M�խ���E܃}� u3��   �M���}���E�    �E�P������躁���E�������Qhĥ �M������E� �������:���jh'  �M�耊���E�E�j hH������赍���E�������P�M������E� ����������ǅ����   �E������M��Ҁ��������R��P���؃��XZ�M�d�    Y_^[�M�3�躥����D  ;��@�����]� ��   �����   �main �����������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q�B`�Ѓ�;�������EPj��MQ�U�R��c�H�Qd�҃�;��X����E�_^[���   ;��E�����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q�Bl�Ѓ�;��ώ��_^[���   ;�迎����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q@�Bh�Ѓ�;��_���_^[���   ;��O�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP��c���   �M��B|��;�����_^[���   ;��܍����]� ����������������������U��j�h&�d�    P��T  SVWQ�������U   ������Y�XD3�P�E�d�    �M�M�����E��}� u3��w  hĥ �M������Eԃ}� u3��Z  �E�P�M������E�    �E�    ������P�M��貝���������������������E�    ������R�M��,�%����E�����������腗���M��,訖���E�P�M�Q�M��B�������   �M������=�   t�׋M������E��}� u��Q���$h'  �M�計��Q�$h'  �M��,������������Iz��������P�M��������������������������E�   ������R�M��,�ɀ���������E�����������贖����������t�M��,�̕�������   R��P�d�Q��XZ�M�d�    Y_^[��`  ;��Ë����]� �   l����   �����   �����   �id data brw ����������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��j���_^[���   ;�赊����]������������������U����   SVWQ��4����3   ������Y�M��M�莏��_^[���   ;��e�����]������������������U����   SVWQ��4����3   ������Y�M��M��̡��_^[���   ;�������]������������������U����   SVWQ��4����3   ������Y�M��M��w���_^[���   ;��ŉ����]������������������U��j�hh�d�    P���   SVWQ������6   ������Y�XD3�P�E�d�    �M�j�M��9����E�    �M��Ov���E������M��	���R��P��|��XZ�M�d�    Y_^[���   ;�������]Ë�   ����    _Lock ����������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��8 td�E���9�tZ�E���M�E�8 t�E�;M�t�E����M���E�8 uh�   h�h\�������E�M��Q��E��     _^[���   ;��!�����]����������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��֟���E�_^[���   ;�讇����]� ������������������������U����   SVWQ��4����3   ������Y�M��EP�M��ɰ���E��M�Q�P�E�_^[���   ;��B�����]� ����������������������������U����   SVWQ��4����3   ������Y�M��EP�M��y����E�_^[���   ;��ކ����]� ������������������������U����   SVWQ��4����3   ������Y�M��EP�M�讇���E�_^[���   ;��~�����]� ������������������������U��j�h��d�    P���   SVWQ������6   ������Y�XD3�P�E�d�    �M�E�M�;t6j�M��݃���E�    �M���r���E�Q�M��ӄ���E������M�蟮���E�R��P�|�;y��XZ�M�d�    Y_^[���   ;�譅����]� �I    �����   �_Lock ����������������������������������������������������������U��j�hȢd�    P���   SVWQ������6   ������Y�XD3�P�E�d�    �M�E�;MtQj�M��ς���E�    �M���q���} t�E�8�t�E�M��P�E�M��E�M��E������M��v���R��P���x��XZ�M�d�    Y_^[���   ;�臄����]� �   �����   �_Lock ����������������������������������������������������������������������U��j�hW�d�    P��  SVWQ��h�����   ������Y�XD3�P�E�d�    �M�ǅx���    �E�    �E�EԋE�P�ys�����EȋE�Ph'  �M�I�����蛫���M��蛠���E��E�;E���  �E�   �E�E��}� ��  �E�E��M��H����E��}� u3���  �M�����E��}� u3��  hĥ �M���}���E��}� u3��  �M���m���Eԉ�t�����t����{����t����E�;E���  �EPj*�M��L�����x���P�M���y�����p�����p�����l����E�    ��l���R�M�� �֚���E�������x����6�����t��� �`  ������P�M��������p�����p�����l����E�   ��x�������x�����l���P�M�� ��r���ȅ�u&�M�� �z���谠��9�t���uǅh���    �
ǅh���   ��h����������E�������x�����t��x�����������v������������}  ǅh���    ǅ\���    ���\�������\�����\���;E��8  ǅP���    ������P�M��������p�����p�����l����E�   ��l���R�M��,�z����E������������ڋ����M��,袝��������P�M��諑����p�����p�����l����E�   ��l���R�M��,�u���������E������������x�����������t?��\�����Ч �M��,�1y����w���;�tǅP���    �ǅP���   ��V�����P��� t�M���|������t��\���Ч ��h��������j,��������������E�   ������ tO��h���P��t����w������̉�����P������p�����t���Q������������l�����l�����h����
ǅh���    ��h����������E�������������D���Q���$h'  ��D����K������m����D���P�M�� ���ԉ����Q���������p��������P�M��跚����l���������������t����B�����t������t����/�����t����M�� 裛�������M���o���j  �EPj*�M��u�����$���P�M��袍����p�����p�����l����E�   ��l���R�M�� ������E�������$����_�����M�� �'�����D���P�M���0�����p�����p�����l����E�   ��l���R�M�� �s����;����E�������D����������;�������   �M�� �v����Ȝ��9�t���t[�M�� �v����������苐���E�� ���̉�X���P�?�����p�����d���Q�M���Ś����l�����d����{������t��� t��t���赒����t���������M��]n���E�    �EȉE��}u�EP�M��:w���EP�MQ�UR�M���m��R��P����p��XZ�M�d�    Y_^[�Ę  ;��N}����]�    �D���   �lodData ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q�B`�Ѓ�;��{����E�P�MQ��c�B�Hp�у�;���z���E�_^[���   ;���z����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���c���   ��M��BT��;��z��_^[���   ;��qz����]������������������������������U����   SVWQ��4����3   ������Y�M���c���   ��M��Bx��;��z��_^[���   ;��z����]������������������������������U����   SVWQ��4����3   ������Y�M���c���   ��M��B(��;��y��_^[���   ;��y����]������������������������������U����   SVWQ��4����3   ������Y�M���c���   ��M��B4��;��1y��_^[���   ;��!y����]������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��Ǡ���E��M�Q�P�E�_^[���   ;��x����]� ����������������������������U����   SVWQ��4����3   ������Y�M��EP�M��e����E�_^[���   ;��Nx����]� ������������������������U����   SVWQ��4����3   ������Y�M��EP�M��Vi���E�_^[���   ;���w����]� ������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �EP�M��x���E�_^[���   ;��{w����]� �������������������������������������U��j�hy�d�    P���  SVWQ��������   ������Y�XD3ŉE�P�E�d�    �M荅���P�M��莇������������������E�    �����R�M�� �����E�����������a�����D���P�M���?�������������������E�   �����R��0���P�M���#����� ����� ����������E���������j����'����E���0��������E�������D����Հ����'�����t�M�� ������X���P�M��賄������������������E�   �����R�M��,�����E�������X����p����M���P�M�'�����u3���  �M�v`���E܋M�>����EЃ}� u3���  hĥ �M��*p���Eă}� u3��  �M�N����E��E�    �E�    �M��b���E�   ��h�����a���E�ǅ\���    ���\�������\����M������9�\���s��\���Ч P�M��i����ȋM���q�������0  ��l���P�M���a�������������������E������R�M��,�׌���E���l����:���M��,�]~���M��,��l����E���=Ч ��   �M��,��l��������P�������e���E�������P�M��,�l��������P�M��Nw���E��������v���������P�M��賂������������������E������R�M��,�md���������E��������p~����������t��M��,�}���$����E�P��L����|i��ǅ@���    ǅ4���    ������P�M���$�������������������E�	�����R�M��,脋���E���������}����M��,诏��������P�M��踃������������������E�
�����R�M��,�g���������E��������}������������  �E�P��$����h����@���P��4���Q��$����,s����t�M��,� k����f���9�4���u��ŋ�@�����y��=�   t�6�����@�����g������������ u����j j��4���P�������Ճ��Pj jh'  �����������P������J����E��}� tj �E�P�����貈������  �}� ��   �E�   j�����P�]��������������������E������R��h����ϑ���E��������a��jj��h���萙��jj��h����7k��j j
��h����r���j j��h����k��j hL��(����Tn���E���(���Pj��h���������E���(���螉��j hL��@����n���E���@���Pj��h����ň���E���@����e���h"  ��t�������P��d����1����E���d���P��h���Q�����R�M�����������[����E���d����ə����[�����tBǅ����    �E������襙���E���h�����`���E������M��`���������  j j��4���P�������΁��Pj jh'  ������蹁��P�������C�������������������E������R������y����E������������}� tj �E�P������x�������  �}� ��   �E�   j������P��Z��������������������E������R�M�蘏���E���������_��h)D j�M��Y���Q���$j�M��3]��Q�H�$j�M��]��Q���$j	�M��]��htemfj�M�����jj
�M��
���j j�M��h��������P�M��,�qg���舀������������������E������Rj�M�胆���E��������#���h"  �����袎��P����������E������P�M�Q�����R�M�ς�������������E������芗���������t?ǅ0���    �E�������f����E���h����^���E������M��r^����0����_�E�������1���������E����U�
�EP�MQ�UR�M��'l����<����E���h���� ^���E������M��^����<���R��P��)�a��XZ�M�d�    Y_^[�M�3��������  ;��m����]� �   �)����   *h���   *L���   *@���   *4���   *$���   *���   *cid brw id data brw bc3 bc2 ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���c���   ��M��B��;��!j��_^[���   ;��j����]������������������������������U����   SVWQ��4����3   ������Y�M��E��M��E��@    �E��@    �E�_^[��]� ���������������������U����   SVWQ��4����3   ������Y�M��E��M��E��M�H�E��M�H�E�_^[��]� �����������������������U���   SVWQ�� ����@   ������Y�M��E�    �EP�M�_����uj�M��]����uǅ ���    �
ǅ ���   �� ����M��}� u�EP�M�l���,  j j ��j�����E�}� u
��   ��   �M�ވ��P�M���u���M������E�jh�'  �M��b��Q���$h'  �M��������pd��Q�$h'  �M��"V��Q���$h'  �M�̄�����Ed��Q�$h'  �M���U��Q���$h'  �M衄�����d��Q�$h'  �M���U��hĥ �M�|������~b���EȋE�Phĥ �M��a������Y���E��-�}� t��E�P��c�Q@�BH�Ѓ�;��g���E�    3�_^[��   ;��vg����]� ����������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH���   �у�;��f��_^[���   ;��f����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH���   �у�;��8f��_^[���   ;��(f����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH���   �у�;��e��_^[���   ;��e����]� ����������������������������������U��j�h��d�    P���   SVWQ������;   ������Y�XD3�P�E�d�    �M��E�    j �M��d��� ����������'  t�}j�M�d��� P�MQ��   ���E��}� u3��oQ���$h'  �M�� a��Q�$������;g���E�    �����P�M�JQ���E�����������r���E����U�
�EP�MQ�UR�EP�M���V���M�d�    Y_^[���   ;��gd����]� ���������������������������������������������������������������������������������U����   SVW��(����6   ������M茀���E��}� u3��=hĥ �M��{^���E�}� u3��#�EP�M��*i��=�   t3���EP�M��K^��_^[���   ;��c����]���������������������������������������������U��j�hF�d�    P��  SVWQ�������E   ������Y�XD3�P�E�d�    �M��E�    j �M�b��� ������������'  t�J  j�M�b��� P�MQ��������E��}� u3��9  �M�P���Q�$h'  �M��P���E����U�
������P�M���>q���������������������E�    ������R�M�� �z���E�������������l����M�� ��~�������P�M����r���������������������E�   ������R�M�� �V��������E�����������l���������t?�M�� �^Z����q����j�M�ba��;0u�E�P�M�� �8Z����i^����V����EP�MQ�UR�EP�M��U���M�d�    Y_^[��   ;��wa����]� ���������������������������������������������������������������������������������������������������������������������������������U���  SVWQ��h����f   ������Y�M��M�g}���E�}� u3��  j h'  �M��,]�����~  hĥ �M��<[���E��}� u3��f  �E�    �EP�,P�����E�3ɋEȺ   �������Q�������l�����l����E��E�P�M��V���E�    �E�P�M�Q�M��`����tK�M��Ug��=�   t�ۋM��oU���E��}� u��Q���$h'  �M��\���EԋM����Eԃ��E��ǅ|���    ���|�������|�����|���;E�}p��D���P�M�|����|����M���ٝP�����|����M���ٝ`�����D���P�M訁����ٝ`�����|����M���ٝd�����D���P�M�����v����E���x�����x���Q�:u�����   R��P�,8�}R��XZ_^[�Ę  ;���^����]�    48����   o8����   j8����   g8D���0   d8ml id data brw �������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�Bp�H\�у�;���]��_^[���   ;��]����]� �������������������������������������U���  SVWQ�������A   ������Y�M���E�P�� ���Q��c�BH�H@�у�;��H]���   ���}�E_^[��  ;��)]����]� �����������������������������������U����   SVW��4����3   �������E�    �M��T���E�} t�M�q���E�E����E���E�_^[���   ;��\����]������������������������������U��j�h��d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M�E�� T�E�   �M��,��f���E��M�� �f���E� �M���VG���E������M��@S���M�d�    Y_^[���   ;���[����]��������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��N��_^[���   ;��e[����]������������������U����   SVWQ��4����3   ������Y�M��M���{��_^[���   ;��[����]������������������U����   SVWQ��4����3   ������Y�M��M��^���E��t�E�P�]N�����E�_^[���   ;��Z����]� ������������������������U��j�h�d�    P���   SVWQ������6   ������Y�XD3�P�E�d�    �M��E�    �M����F���E��M���kb���E��E�M��EP�M���Qu���E�M�H(�E������M�ir���E�R��P�\=�YM��XZ�M�d�    Y_^[���   ;���Y����]� �   d=����   p=_$ArrayPad ���������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ��c�B�Hp�у�;��Y���E�_^[���   ;��Y����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q�B`�Ѓ�;��X���E�_^[���   ;��X����]�������������������������U��j�h+�d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M��E�    �M���p���E������M���`H���M�d�    Y_^[���   ;���W����]��������������������������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �E���P�M�d����,�������,����E_^[���   ;���V����]� ����������������������������U����   SVWQ��4����3   ������Y�M��E��@(_^[��]�����������������U����   SVWQ��4����3   ������Y�M��EP�M����jv��_^[���   ;��>V����]� ������������������������U��j�h��d�    P��l  SVW��������   ������XD3ŉE�P�E�d�    �M��W���E�E�P�M�e���E�    �E�P�tE�����E��E�    �E�    ��h0 �|@��P�M���Q��c�B��H  �у�;��sU���E���h0 �|@��Pj��c�Q��H  �Ѓ�;��CU���E��M���q���E�Q���$h'  �M��DQ���E��XQ���$h'  �M��+Q���E��XQ���$h'  �M��Q���E��hĥ �M��O���E��E�P�M��J��ǅx���    �Eă���`�����x���P��l���Q�M�� U����tk��x�����[��=�   t�ҋ�x�����I����T�����T��� u�Q���$h'  ��T����{P���Zv����`����U�����`�������`����{���j h( ������� Q���E�j h  �������
Q���E����􉥘���������P�M�Q������R������P��h�����������������������E�������RV��h�����������M�\O���E��������l���E���������k���E� ��������k�����̉�����j h �bP���������M�
O��ǅH���    ���H�������H�����H�����   �M�o��j h ������P���E��������������Pj0j j�j���H����U�Q���$�����P�h�����������������������E�������RV�g�����������M�WN���E�������k���E� �������j���6������̉�4���j h �gO���������M�N�����̉�@���j h  �BO���������M��M��ǅ<���    ���<�������<����Eă�9�<���}w�M�zn�����ĉ�L�����<����U���QP��r�����������M�M���Eă�9�<���t-�M�5n�����̉�X���j h��N���������M�OM���l����M�n�����̉�d���j h��uN���������M�M�����̉�p���j h��PN���������M��L���E������M��i��R��P�(F�D��XZ�M�d�    Y_^[�M�3��yf����x  ;���P����]ÍI    0F����   lF����   hFx���   cFl���   `Fid data brw knotennameC4D ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h
�d�    P���   SVW������;   ������XD3�P�E�d�    ǅ,���    �EP�MQ�������[������������������E�   �������_��P�M�[����,�������,����E� ������
g���E�M�d�    Y_^[���   ;��}N����]����������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M���_��P�M��yi���E�_^[���   ;���M����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q�B�Ѓ�;��M��_^[���   ;��M����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H�Q0�҃�;��M��_^[���   ;��M����]� ����������������������������������U����   SVW��$����7   ��������̉�,���j h� �I����$����M�QH�����̉�8���j h� �I����$����M�,H��_^[���   ;��hL����]�������������������������������������U��j�hS�d�    P��8  SVW�������N   ������XD3ŉE�P�E�d�    j h� �M���H���E�    �M��MY����u$ǅ����   �E������M��4d���������   j h� �������H���E�j ���̉�����j h� �H��������������PhϦj�M�Qhå �s����(�������������������E� �������c�������� t!ǅ���   �E������M��c��������ǅ���    �E������M��qc�������R��P�`L�^>��XZ�M�d�    Y_^[�M�3��@`����D  ;���J����]Ë�   hL����   tLname �������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M���[�������_^[���   ;���I����]����������������������������U����   SVW��0����4   ������h� j+hij8�wT������8�����8��� t��8����O����0����
ǅ0���    ��0���_^[���   ;��jI����]���������������������������������������U��j�h��d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M�M��d���E�    �E�� T�M���*6���E��M�� ��P���E��M��,��P���E������E�M�d�    Y_^[���   ;��H����]�����������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��'L���E�� 4!�E�_^[���   ;��H����]����������������������U����   SVWQ��4����3   ������Y�M��M��?���E��t�E�P�];�����E�_^[���   ;��G����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��`���E�� �!�E�_^[���   ;��IG����]����������������������U����   SVWQ��4����3   ������Y�M��M��9���E��t�E�P�:�����E�_^[���   ;���F����]� ������������������������U����   SVW�� ����8   ������} w	�E    �+���3��u��sj ��$����]��h<���$���P�k��jVh("�l��P�EP�h5������8�����8���_^[���   ;��3F����]������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M���L���E�� �"�E�_^[���   ;��E����]� �������������������������������U����   SVWQ��4����3   ������Y�M��E�� �"�M���V��_^[���   ;��LE����]�������������������������U����   SVWQ��4����3   ������Y�M��M���4���E��t�E�P�8�����E�_^[���   ;���D����]� ������������������������U����   SVWQ������;   ������Y�M��} w	�E    �+���3��u��sj ������[��h<������P�i��jah("�j��P�EP�c3������,�����,���_^[���   ;��.D����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��EP�W����_^[���   ;���C����]� ���������������������������U��j�h�d�    P���   SVWQ������6   ������Y�XD3�P�E�d�    �M�Q�̉� �����.���M��]���E�    �M��X���M�A�E��@    �E������E�M�d�    Y_^[���   ;��C����]�������������������������������������������������U��j�h�d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M��E�    �M��$H���E������M��>`���M�d�    Y_^[���   ;��UB����]����������������������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �E�P�M��QR�Z����� P�M�>����,�������,����E_^[���   ;���A����]� �����������������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �E�P�M��QR�M�>����,�������,����E_^[���   ;��>A����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E�3Ƀx ����_^[��]�������������������������U��j�hg�d�    P���   SVWQ�������>   ������Y�XD3�P�E�d�    �M�ǅ ���    �E�   �EP���̉�����UR�UU���� ����M��H@���M��E�����̉����P�.U���� ����EP�M��HL���������� ������� ����E� �M�`Y���E�M�d�    Y_^[��  ;��?����]� �����������������������������������������������������������������������U��j�hҨd�    P��  SVWQ�������C   ������Y�XD3�P�E�d�    �M�ǅ���    �E�   �E;E�u�E�M;Huh  h�"h�"�X����j ������P�M�H���������������������E��������5���E��E��������4X���E�P�M�Q�M��3���E�M�;H��   �E�P��V�������M�Q��:�����R��V�������E�P��:�������M�Q��V�����R�:�������E�P�M����h��j�E�P�M���7F���E�H���U�J���̉�����EP�S���������MQ�M��5J���������������������E� �M�MW���E�M�d�    Y_^[��  ;��=����]� ��������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M�� '���E�_^[���   ;���<����]�������������������������������U����   SVWQ��4����3   ������Y�M��M��_��_^[���   ;��u<����]������������������U����   SVWQ��4����3   ������Y�M��M���N���E�_^[���   ;��"<����]�������������������������������U����   SVWQ��4����3   ������Y�M��M���A���E�_^[���   ;���;����]�������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��~[���E��M�P3�;Q��_^[���   ;��P;����]� ��������������������������U����   SVWQ��4����3   ������Y�M��EP�M��+���������_^[���   ;���:����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��EP�M���F���E�� �"�E�_^[���   ;��u:����]� �������������������������������U����   SVWQ��4����3   ������Y�M��M��\I���E�_^[���   ;��:����]�������������������������������U����   SVWQ��4����3   ������Y�M��M��P��_^[���   ;��9����]������������������U����   SVWQ��4����3   ������Y�M��M��.��_^[���   ;��e9����]������������������U����   SVWQ��4����3   ������Y�M��M���>��_^[���   ;��9����]������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��@����0   ������E��_^[��]����������������������U��j�h7�d�    P���   SVWQ������6   ������Y�XD3�P�E�d�    �M�ǅ ���    �E�   �E�P�MQ�M�4���� ������� ����E� �M�gQ���E�M�d�    Y_^[���   ;��7����]� ����������������������������������������������U��j�hx�d�    P���   SVWQ������9   ������Y�XD3�P�E�d�    �M��E�    �E;E�th�  h�"h�#�BP�����M��-���E��EP�M�Q�3�����R�E�P�M��;*���E�j�M��C3���E�P�X3�����Mԉ�E�P�G3�����Q�CO�����Uԉ�E������M�:P���M�d�    Y_^[���   ;��z6����]� ��������������������������������������������������������������������U��j�h��d�    PQ���   SVWQ������:   ������Y�XD3�P�E�d�    �e��M�j�M����B���E��E�    �E�    �E�P�ZN����������M�Q�����R�M���:���EЃ��EЋE�P�"2����������M�Q�����R�M���:���E�}� ~�E�P��M����P�M���LU��j�E�P�M���{=��j j �xZ���E�������a��E������E�R��P�0b�(��XZ�M�d�    Y_^[���   ;���4����]Ë�   8b����   Db_Pnode �����������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��C;���E��HQ��L����P�M����#T���E��HQ�0����P�M����T��j�E��HQ�M����4<���E��@    _^[���   ;���3����]����������������������������������������������U����   SVWQ������9   ������Y�M�j�M��X1���E�E��E��8 tJ�E���U��A;Bt�} t�E���Q;Ut�E�����M���E���    �E���U��A�뮍M���[��R��P�$d�&��XZ_^[���   ;��3����]�    ,d����   8d_Lock ������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M�Q�̉�,����EP��X���M��XQ���EP�M�����X���E�_^[���   ;��A2����]� ���������������������������U����   SVWQ��4����3   ������Y�M��M���@��_^[���   ;���1����]������������������U����   SVWQ��4����3   ������Y�M��M��2��_^[���   ;��1����]������������������U����   SVWQ������9   ������Y�M�j�M��(/���E��8�t3�E��E���E���U��A��E��8 t�E���    �ދE��     �M���Y��R��P�8f�r$��XZ_^[���   ;���0����]ÍI    @f����   Lf_Lock ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVWQ��4����3   ������Y�M��EP��#����_^[���   ;��!0����]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�$:����_^[���   ;���/����]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M��M6���E�_^[���   ;��Z/����]� ��������������������U����   SVWQ��4����3   ������Y�M��M��y���E��@    �E�_^[���   ;���.����]���������������������U����   SVWQ��4����3   ������Y�M��E��8 t�E��x t�E���U��B;Auch�   h�"hX%�G�����   ��tC3�u!h�$j h�   h�"j�K ������u�j h�   h�"h $h�#�14�����E��HQ��Q����_^[���   ;��.����]�������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 t�E��x t�E���U��B;Auch�   h�"h�&�F�����   ��tC3�u!h�$j h�   h�"j�K������u�j h�   h�"h�%h�#�13�����E��HQ��E�����U�� �B�E�_^[���   ;��-����]������������������������������������������������������������U��j�h��d�    P���   SVWQ������;   ������Y�XD3�P�E�d�    �M�ǅ���    �E�P�M��A���E�   �M���>���E�P�M�A���������������E� �M���E���ER��P�k���XZ�M�d�    Y_^[���   ;��,����]� �   k����   (k_Tmp �������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 t0�E��x t'�E��HQ� (�����U�� �B�M���E��H;Juch  h�"h�'�xD�����   ��tC3�u!h�$j h  h�"j�������u�j h  h�"h�&h�#��0�����E�_^[���   ;���*����]������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��8 t�E��M�;tch<  h�"h�)�LC�����   ��tC3�u!h@)j h=  h�"j��������u�j h=  h�"hX(h$(�/����_^[���   ;��)����]� ������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��
>���E�_^[���   ;��>)����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��R���E�_^[���   ;���(����]�������������������������������U����   SVWQ��4����3   ������Y�M��M��B���E�_^[���   ;��(����]�������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E�_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVW��@����0   ������E��_^[��]����������������������U����   SVWQ������9   ������Y�M�j �E�P�M�����E��HQ��?������U��E��HQ��?�����U��J��E��HQ�#�����U��J��E��@    ��E�E��E��M�;Ht3�E�P�?������M�E�P�M����Q��j�E�P�M����/���_^[���   ;��&����]����������������������������������������������������������U��j�h0�d�    PQ���   SVWQ������:   ������Y�XD3�P�E�d�    �e��M�j�M���3���E��E�    �E�    �E�P�>����������MQ�����R�M���+���EЃ��EЋE�P�r"����������MQ�����R�M����*���EЃ��EЋE�P�I����������MQ�����R�M���",���c�}�~�E�P�"����P�M���kE���}� ~�E�P��=����P�M���ME��j�E�P�M���|-��j j �yJ���E�������q��E������E܋M�d�    Y_^[���   ;��%����]� ��������������������������������������������������������������������������������������������������U��j�hk�d�    P��(  SVWQ�������J   ������Y�XD3�P�E�d�    �M�M���A���M�+A;EsLh�)������/���E�    �����P�������7��h��������Q�PI���E������������"���E�HM�U�J�M�d�    Y_^[��4  ;���#����]� ���������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��:���E�� *�E�_^[���   ;��E#����]� �������������������������������U��j�h��d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M�M�� ���E�    �E�� *�EP�M����+���E������E�M�d�    Y_^[���   ;��"����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M������_^[���   ;��""����]�������������������������������U����   SVWQ��4����3   ������Y�M��M��C6���E��t�E�P�]�����E�_^[���   ;��!����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� *�M����K ���M���2��_^[���   ;��A!����]������������������������������U����   SVWQ��4����3   ������Y�M��E�� *�M��Z5��_^[���   ;��� ����]�������������������������U����   SVWQ��4����3   ������Y�M��M�����E��t�E�P������E�_^[���   ;��n ����]� ������������������������U��j�hتd�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M�EP�M��<,���E�    �E�� *�E��P�M���')���E������E�M�d�    Y_^[���   ;������]� �����������������������������������������������������U��j�h�d�    P���   SVWQ������6   ������Y�XD3�P�E�d�    �M�Q�̉� ����g.���M��nB���E�    j j �M��rD���EP�M��	���E������E�M�d�    Y_^[���   ;�������]� ����������������������������������������������U��j�h8�d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M�EP�M��=���E�    j j �M��C���(*Pj �MQ�M���H���E������E�M�d�    Y_^[���   ;������]� ������������������������������������������������U��j�hh�d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M��E�    j j�M���B���E������M��(D���M�d�    Y_^[���   ;��a����]����������������������������������������������U����   SVWQ��4����3   ������Y�M��M��#��_^[���   ;�������]������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;������]������������������U����   SVWQ��4����3   ������Y�M��M��B+��_^[���   ;��U����]������������������U����   SVWQ��(����6   ������Y�M��M�=!��;Es�G���M�+!��+E�E�E;E�s�E�E�E�;Eu%�(*P�MM�Q�M��v;���URj �M��h;���Ij �E�P�M�����ȅ�t4�E�P�M�O"��EP�M��QR�M��94��P�+�����E�P�M������E�_^[���   ;��f����]� ����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M�h<  h0*�EP�q�����EP�w7����P�MQ�M���5��_^[���   ;��~����]� ����������������������������������������U����   SVW��@����0   ������EP��8����_^[���   ;������]�������������������U����   SVWQ��(����6   ������Y�M��E��u�J�E��xrA�E��H�M�} v�EP�M�Qj�U���R�)�����E��H��Q�U�R�M����U*���E��@   �EP�M�����_^[���   ;��c����]� ���������������������������������������������U����   SVWQ��0����4   ������Y�M��E��xr�M��Q��0�����E�����0�����0���_^[��]������������������������������U����   SVWQ��4����3   ������Y�M��M���+���EP�M����?-���E�_^[���   ;��s����]� �����������������������������U����   SVWQ��4����3   ������Y�M��M��b+���E��P�M�����,���E�8�u	�E�� �����E�_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M��M���%���E�_^[���   ;������]�������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��} th,  h0*�EP�	�����EP�M������ȅ�t �EP�M��m/���M+�Q�U�R�M��qA���Dj �EP�M��o���ȅ�t,�EP�MQ�U��BP�M��-/��P�&�����EP�M������E�_^[���   ;��Z����]� ����������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��H;Ms�)���E��H+M;Ms�E��H+M�M�} vR�E��H+M+MQ�M��c.��EEP�U��B+EP�M��J.��EP�,�����E��H+M�M�E�P�M������E�_^[���   ;��h����]� ��������������������������������������������������U����   SVWQ��(����6   ������Y�M�ƅ/��� �E��M�H��/���R�M��-��EP�1����_^[���   ;�������]� ����������������������������U����   SVW��@����0   ������E�M��_^[��]������������������U����   SVWQ��0����4   ������Y�M��M��'��;Es�*4���E��H;Ms�E��HQ�UR�M��17���S�E��t;�}s5�E��M;Hs�U��0�����E��H��0�����0���Rj�M��79����} u
j �M��"��3�;E���_^[���   ;������]� ���������������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��xr�M��Q��0�����E�����0�����0���_^[��]������������������������������U����   SVWQ��4����3   ������Y�M��EP�m����_^[���   ;�������]� ���������������������������U����   SVWQ��(����6   ������Y�M�Q�̉�,����EP��8���M��\���EP�M�����<���E�_^[���   ;��A����]� ���������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVWQ��4����3   ������Y�M�j �EP������_^[���   ;������]� �������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�(����_^[���   ;��=����]� �����������������������U����   SVWQ��4����3   ������Y�M��EP�w����_^[���   ;�������]� ���������������������������U��j�h��d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M�M�������E�    �E�M�H�EP�M��B���E������E�M�d�    Y_^[���   ;��5����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M���.���E�� *�E�_^[���   ;������]� �������������������������������U����   SVWQ��$����7   ������Y�M��M����|���E�}�wǅ$���   ��E����$�����$���_^[���   ;��+����]����������������������������������������U��j�h��d�    PQ���   SVWQ������:   ������Y�XD3�P�E�d�    �e��M�E���E܋M����;E�s�E�E��C�E�H��E�3Ҿ   ��;�s+�E�p��M��V��+ƋM�9Aw�E�H��U�J�M��E�    �E�    �E܃�P�M������������������M��f�e��E�E��E��E܃�P�M�����������������M��"j j�M��I3��j j �"3���E�   �Q���E�   �E�   �e���E������} v �EP�M��T&��P�M܃�Q�U�R�����j j�M���2���E�MЉH�E�M܉H�EP�M������M�d�    Y_^[���   ;��P����]� ��������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��} t �M��J%��9Er�M��=%���M�A;Ew2����_^[���   ;��o����]� �������������������������U����   SVWQ��4����3   ������Y�M��M������_^[���   ;������]�������������������������������U����   SVWQ��(����6   ������Y�M�Q�̉�,����EP�52���M��,���EP�M�����1���E�_^[���   ;������]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ��.����_^[���   ;��-����]� �����������������������U����   SVWQ��4����3   ������Y�M�j �EP�4����_^[���   ;���
����]� �������������������������U����   SVWQ��$����7   ������Y�M��E������}� v�E쉅$����
ǅ$���   ��$���_^[��]�������������������������������U����   SVWQ��4����3   ������Y�M��M��9���E�_^[���   ;��
����]� ����������������������������U����   SVWQ��$����7   ������Y�M��E����?�}� v�E쉅$����
ǅ$���   ��$���_^[��]�������������������������������U����   SVW��@����0   ������} u�EP�MQh�*�q"����_^[���   ;��'	����]��������������������U����   SVW��@����0   ������} t�EP������_^[���   ;�������]�����������������������������U����   SVW��4����3   �������Q����;�����;���P�MQ�UR�EP�MQ�����_^[���   ;��W����]������������������������������������U����   SVW��@����0   ������_^[��]������������U����   SVW��4����3   �����������;�����;���P�MQ�UR�EP�MQ�����_^[���   ;������]������������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVW��,����5   ������} w	�E    �+���3��u��sj ��0������h<���0���P�',���Ek�P�����_^[���   ;�������]��������������������������������������U����   SVW��$����7   ������E�E��E�Pj��������,�����,��� t��,����U����,�����$����
ǅ$���    _^[���   ;��*����]���������������������������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��@����0   ������_^[��]������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVW��$����7   ������E�E��E�Pj�������,�����,��� t��,����U����,�����$����
ǅ$���    _^[���   ;�������]���������������������������������������U����   SVW��,����5   ������} w	�E    �+���3��u��sj ��0�������h<���0���P�)���EP������_^[���   ;��<����]�����������������������������������������U����   SVW��4����3   ������E�R��P�L��Q���XZ_^[��]ÍI    T�����   `�_Secure ������������������������U����   SVW��@����0   ������EP�MQ�UR�EP��+����_^[���   ;��Z����]�����������������������U����   SVW��@����0   ������EP�MQ�UR�EP� �����E_^[���   ;�������]��������������������U����   SVW��@����0   ������EP�MQ�UR�EP�����_^[���   ;������]�����������������������U����   SVW��@����0   ������EP�MQ�UR�EP��"�����E_^[���   ;��7����]��������������������U��j�h�d�    P��,  SVWQ�������K   ������Y�XD3ŉE�P�E�d�    �M�M�u���E܃}� u3��y  �E�E�j h4+�����������E�    ������P�M������E����������������E�P�������E�   jj�M��_)��jj�M��	���Q���$j�M��-���Q���$j�M�����Q���$j�M�����Q���$j �M������j h'  �M���)��Ph'  �M���(��j h'  �M���)��������������
�p  �������$�,�Q���$j�M������N  Q�0+�$Q�,+�$�  ���$j�M��s����   Q���$j�M��^����  Q�(+�$Q�,+�$�k  ���$j�M��0�����   Q�$+�$Q�,+�$�=  ���$j�M������   Q� +�$Q�,+�$�  ���$j�M�������   Q�+�$Q�,+�$��  ���$j�M������VQ�+�$j�M������@Q�+�$j�M��z����*Q�+�$j�M��d����Q�+�$j�M��N���ǅ����   �E������M�����������R��P������XZ�M�d�    Y_^[�M�3������8  ;�������]� ��   �����   (�wc �T�i�����ږ�6�a�w�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������Q�E�$Q�E�$�{�����_^[���   ;�������]�������������������������U����   SVW��<����1   �������E���$�E���$�&����ٝ<���م<���_^[���   ;��<�����]�������������������������U����   SVWQ��$����7   ������Y�M��M����E�} u3��  j h'  �M���%����$�����$���
�p  ��$����$��Q���$j�M������N  Q�0+�$Q�,+�$�������$j�M��]����   Q���$j�M��H����  Q�(+�$Q�,+�$�U������$j�M�������   Q�$+�$Q�,+�$�'������$j�M�������   Q� +�$Q�,+�$��������$j�M������   Q�+�$Q�,+�$��������$j�M������VQ�+�$j�M��z����@Q�+�$j�M��d����*Q�+�$j�M��N����Q�+�$j�M��8����   _^[���   ;��>�����]� j������L�w���������������������������������������������������������������������������������������������������������������������������������������������������U���   SVWQ�� ����@   ������Y�M��E�    �EP�M������uj�M�.�����uǅ ���    �
ǅ ���   �� ����M��}� u�EP�M������  j j �)������E�}� u
�>  �9  �M��}���EԋM�r���EȋM���P�M�����jh�'  �M��^���j h'  �M��"��Ph'  �M��!��j j�M��y"��Pj�M��t!��j h'  �M��_"��Ph'  �M��W!��j j�M������Pj�M������Q���$j�M��W���Q�$j�M�����Q���$j�M��9���Q�$j�M������Q���$j�M�����Q�$j�M������Q���$j�M������Q�$j�M�����Q���$j �M������Q�$j �M������E��-�}� t��E�P��c�Q@�BH�Ѓ�;������E�    3�_^[��   ;��m�����]� ���������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P��  SVW��8����/  ������XD3ŉE�P�E�d�    �M�������3���E�M�������E�    j j�M�������Eă}� tHj h�+�������V�����x�����x�����t����E���t���Q�M��r���E� ����������Fj h�+������������x�����x�����t����E���t���Q�M��*���E� �������K���M������E�j j�M������x�����x�������x�����x����|  ��x����$�h�j h�+������������x�����x�����t����E���t���Q�M�����E�����������$  j h�+�������6�����x�����x�����t����E���t���Q�M��R���E��������s����   j h�+�������������x�����x�����t����E���t���Q�M�����E��������(���   j h�+������������x�����x�����t����E���t���Q�M�����E������������Fj h�+������X�����x�����x�����t����E���t���Q�M��t���E������������̉�(���j h�+������x����M�����M���j h� ��@���������E�	j h�+��p���������E�
j h�+�����������E�j h�+�����������E�����4�����@���Pj0j j�j�Q���$j�M�����Q�$��X���Q�
������x�����x�����t����E���t���P��p���Qj0j j�j�Q���$j�M��J���Q�$������R��	������p�����p�����l����E���l���Q������Rj0j j�j�Q���$j�M������Q�$������P�	������h�����h�����d����E���d���R������P������Q�������`�����`�����\����E���\���P�� ���Q�s������X�����X�����T����E���T���P�����Q�G������P�����P�����L����E���L���P��0���Q�������H�����H�����D����E���D���P��H���Q��������@�����@�����<����E���<���PV��������8����M�c����E���H�������E���0���� ���E��������
���E��� �����
���E���������
���E���������
���E��������
���E���X����
���E��������
���E�
�������
���E�	��p����y
���E���@����j
��j h ��l���������E�j h|+������������E�����`�����l���P�M�Q������R������P�������x�����x�����t����E���t���RV�������p����M�#����E���������	���E���������	���E���l����	��j h �������.����E�j ht+�����������E����􉥴���������Pj0j j�j�Q���$j�M�����Q�$������Q�������x�����x�����t����E���t���P������Q�����R�������p�����p�����l����E���l���QV�������h����M�&����E�����������E������������E�����������E����������j hp+��,����"����E�j hd+��D��������E����� �����,���P�M�Q��D���R��\���P��������x�����x�����t����E���t���RV��������p����M�^����E���\����
���E���D��������E���,�������j h �������i����E�j hP+�������S����E� ����t���������Pj0j j�j�Q���$j �M��I���Q�$������Q��������x�����x�����t����E�!��t���P������Q������R��������p�����p�����l����E�"��l���QV��������h����M�a����E�!����������E� �����������E������������E������������M�������̉�����j h� �P�����x����M������E� �M�����E������M����R��P�4�����XZ�M�d�    Y_^[�M�3��m�����  ;��������]ÍI    <�����   [�����   T�type_S headlight_S ���֠!�l���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E�� �+�M��&���_^[���   ;��������]�������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�������E�_^[���   ;��^�����]� ������������������������U��j�hc�d�    P��8  SVW�������N   ������XD3ŉE�P�E�d�    j h�,�M�������E�    �M��M�����u$ǅ����   �E������M��4���������   j h�,�����������E�j ���̉�����j h�,����������������Ph�j�M�Qh¥ �����(�������������������E� ��������������� t!ǅ���   �E������M����������ǅ���    �E������M��q�������R��P�`��^���XZ�M�d�    Y_^[�M�3��@�����D  ;��������]Ë�   h�����   t�name �������������������������������������������������������������������������������������������������������U����   SVW��0����4   ������h�,jhij���������8�����8��� t��8����	�����0����
ǅ0���    ��0���_^[���   ;��������]���������������������������������������U����   SVWQ��4����3   ������Y�M��M�����E�� �+�E�_^[���   ;��Y�����]����������������������U��j�h��d�    P��\  SVWQ��������   ������Y�XD3ŉE�P�E�d�    �M�E��u3��_  �M��
����E�    jdh�   j�j��M��.������  �E�P�MQ�UR�������=����E�������������t�������M����u3ǅ���������E� �������c����E������M�������������  h1D4ChCD4Cjj j�EP�������������q�����uA�����������������������E� ������������E������M������������^  ���������������������������������������t������P������������P�MQ����������̉�����j hL�����������������������E�jj�������w�����0�   ����󥍍�����8���������P������Q�E��  ��P������"����������+�����0����t"j jj�M�c���P�EP������Q�E��������������������� ����E� �����������E������M��U����� ����ǅ���    �E������M��4��������R��P�в�����XZ�M�d�    Y_^[�M�3��������h  ;��W�����]� �   ز����@   �������   �vrml startDialog ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���  SVWQ�������G   ������Y�M��M������M��������M���������M���$�����Q���$Q���$Q���$����������M����P�Q�@�AQ���$Q���$Q���$�����������M������P�Q�@�AQ���$Q���$Q���$���������M������P�Q�@�AQ���$Q���$Q���$��$����w���M���$���P�Q�@�A�E�_^[��  ;��(�����]�������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E����X�M����Y�U�����E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��E��E��E��E�X�E��E�X�E�_^[��]� �����������������������U����   SVWQ��4����3   ������Y�M��M�������E�� H-�E�_^[���   ;��������]����������������������U����   SVWQ��4����3   ������Y�M��M������_^[���   ;��u�����]������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�������E�_^[���   ;�������]� ������������������������U��j�hy�d�    P��  SVW��D�����   ������XD3ŉE�P�E�d�    �E�P�w  ���E�P�  ���E؋E�P�@������M��D� ���̉�d���j h�-�h�����\����M�������̉�p���j h�-�C�����\����M�����j h �������#����E�    j h�-�������
����E�����|���������P������Q������R�M��������P�����\�����\�����X����E���X���������T�����T�����P����E���P���R������P������Q��������L�����L�����H����E���H���PV�k�������D����M�����E������������E������������E�������������E� �����������E������������r���j h �����������E�   j h|-��H���������E�������������Pj �M�Q��0���������\�����\�����X����E���X���P��H���Q��`���R��������T�����T�����P����E���P���QV�d�������L����M������E���`��������E���0��������E���H��������E�����������z���j jP�E�P������jjN�E�P��x���Q�M�������\�����\�����X����E�	   ��X����=����E�������x����������̉�����j hx-������\����M�=���j������P�M�^�����\�����\�����X����E�
   ��X�������P�U�R�M�������]����E������������������̉�����j ht-������\����M����R��P�T��k���XZ�M�d�    Y_^[�M�3��M����ļ  ;��������]ÍI    \�����   {�����P   t�header ltime �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������EP������_^[���   ;��F�����]�������������������U����   SVW��@����0   ������EP������_^[���   ;��������]�������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�HP�у�;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q�BT�Ѓ�;�����_^[���   ;�������]� �����������������������������U����   SVW��@����0   ������EP�M���   Q�UR������_^[���   ;�������]���������������������U��j�hj�d�    P��4  SVW��������   ������XD3ŉE�P�E�d�    �E�    �} ��  �E�    �E�    �M��/����E@�EЋED�EċM�X������̉�����P�������������t���P�
������������E�ǅh���    ��t���P��P��������E���@���P�M��@�T����������������������E�������R���̉�������P���P�q��������������Q��������������������������E�������P��,���Q�M��@�&����������������������E������������������E���,��������E������������E���@����������������
  j h�-��l��������E���h���P��T���Q�~������������������������E�������P��l���Q��t���R������P�n������������������������E�������R������P�B������������������������E�	������R��P����M����E��������n����E��������_����E���T����P����E���l����A�����h�������h����	�����P���P��t�����������̉�������t���P����������������Q�#������������������������E�
������P������Q�M��@�����������H����E��������)������̉� ���j h �����������M�����j8������������E������ tn���̉�$����EHP������������������������E����̉�0�����t���R�����������EP�E�������l����������������������
ǅ����    ������������E��������D���ǅ8���    �M������,����M������ ����M�G�����������t
ǅ,���    �M�*������������t
ǅ ���    ��,��� u�� ��� u
ǅ8���   ��,��� u�� ���u�}D t
ǅ8���   ��,���u�}@ t�� ��� u
ǅ8���   ��,���u�}@ t�� ���u�}D t
ǅ8���   ��8��� ��   j h�'  �M��������������t!��D���P�MQ�������E�   �E�   �}� u��D���P�MQ�S�����j h�'  �M������������t��D���P�MQ�w������E�   ��D��������=�  u��D���P�MQ��������D��������=�  u(�}� u"��D���P��0�   �u���MQ�������8�E�   �E�   ��E�    �E�    ���ĉ�<���P��D����߻���������������������E��U�R�E�P��0�   �u����M����P�MQ�E�������P��8��� t8j h�'  �M�������q�����t�EP��������}� u�EP�������M�����E��D�����T�����T�����H�����H��� tj��H����l����������
ǅ����    �E���P���������E� ��t���������"����E������MH����R��P������XZ�M�d�    Y_^[�M�3�������@  ;�������]Ë�   �����0   X�t���   J�P���   <�knotennametmp knotennameC4D mg ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M������_^[���   ;�������]������������������U����   SVWQ��4����3   ������Y�M��M��	���_^[���   ;��E�����]������������������U����   SVWQ��4����3   ������Y�M��M��W����E��t�E�P�������E�_^[���   ;��������]� ������������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;�������]������������������U����   SVWQ��4����3   ������Y�M��M������_^[���   ;��5�����]������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��������]������������������U��j�h��d�    P��  SVW��������  ������XD3�P�E�d�    j h4.��P��������E�    j h  �������f����E�����D�����P���P��h���Q�M�8�����<�����<�����8����E���8���P������Q������R��������4�����4�����0����E���0���QV���������,����M�����E��������<����E���h����-����E� �����������E�������P��������M�Q����E�P�M�������P����M؉M�j h �������h����E�   j h �������O����E�j h ������9����E�j h$.��L����#����E����􉥰���������Pj0j j�j��M�Q��$������R��������<�����<�����8����E���8���Q������Rj0j j�j��E�Q�@�$�����Q�e�������4�����4�����0����E�	��0���P�����Qj0j j�j��U�Q�B�$��4���P� �������,�����,�����(����E�
��(���R��L���P��d���Q�>�������$�����$����� ����E��� ���P��|���Q����������������������E������P������Q�����������������������E������P������Q����������������������E������P������Q������������������ ����E��� ���PV�h������������M�����E������������E������������E������������E���|��������E�
��d����r����E�	��4����c����E�������T����E��������E����E���L����6����E�������'����E������������E����������������E�P�M������������M��M�j h �������j����E�   j h ������Q����E�j h ��H����;����E�j h.��x����%����E���������������Pj0j j�j��M�Q�A�$�� ���R��������<�����<�����8����E���8���Q�����Rj0j j�j��E�Q�@�$��0���Q�f�������4�����4�����0����E���0���P��H���Qj0j j�j��U�Q��$��`���P�"�������,�����,�����(����E���(���R��x���P������Q�@�������$�����$����� ����E��� ���P������Q����������������������E������P������Q�����������������������E������P������Q����������������������E������P������Q������������������ ����E��� ���PV�j������������M�����E������������E������������E������������E������������E��������t����E���`����e����E���0����V����E��� ����G����E���x����8����E���H����)����E�����������E����������������E�P�M�������x�����`����e�����t���P��`���Q�U�R蜰����j h ������M����E�   j h ��D����4����E�j h ��t��������E�j h �����������E�j h.������������E� ������������Pj0j j�j�Qمt����$��,���Q�x�������<�����<�����8����E�!��8���P��D���Qj0j j�j�Qم`����$��\���R�3�������4�����4�����0����E�"��0���Q��t���Rj0j j�j�Qمd����$������P���������,�����,�����(����E�#��(���R������Pj0j j�j�Qمh����$������Q��������$�����$����� ����E�$�� ���P������Q������R�����������������������E�%�����Q�����R����������������������E�&�����Q�����R�o���������������������E�'�����Q��4���R�C����������������� ����E�(�� ���Q��L���R�������������������������E�)������Q��d���R��������������������������E�*������Q��|���R�������������������������E�+������QV�������������M�3����E�*��|���������E�)��d���������E�(��L���������E�'��4��������E�&����������E�%����������E�$�����������E�#�������v����E�"�������g����E�!��\����X����E� ��,����I����E��������:����E��������+����E���t��������E���D��������E����������������M�@������̉�����j h .�k�����<����M�����M����R��P���蹴��XZ�M�d�    Y_^[��  ;��+�����]ÍI    �����   S�����   O�����0   K�t���   E�`���   @�axis angle ml1 $S2 $S1 ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ�� ����8   ������Y�M���E�P��$���Q��c�BH�H(�у�;��x����U��
�H�J�@�B�E_^[���   ;��R�����]� ��������������������������������������������U����   SVWQ�� ����8   ������Y�M���E�P��$���Q��c�BH�H0�у�;��ؼ���U��
�H�J�@�B�E_^[���   ;�貼����]� ��������������������������������������������U���\  SVW�������W   ������u�   �}��E�P������Q���������U؋H�M܋P�U��E�P������Q���������U�H�M�P�U�E�P������Q��������U��H�M�P�U��E��E��E��%X.�5H.���$�������E��E��e�E��E��e��E�X�E��e܋E�X�EP������Q�<������U��
�H�J�@�BQ���$�EP���������t7Q���$Q���$Q���$�������k����M���P�Q�@�A�E���R��P��荮��XZ_^[��\  ;��
�����]Ë�   $�����0   0�m ��������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ���������]����Az���+��x.�]����u�h.����E�$蛼����_^[���   ;�������]������������������������������������U����   SVW��(����6   ������E� �M�	�U�B�E�H���M�A�U�J��ٝ0���م0���Q�$�N������]��E���.����DzQ���$�M�����E�_�E������]��E�@�M�ٝ0���م0���Q�$�M�A�M�ٝ,���م,���Q�$�U��M�ٝ(���م(���Q�$�M�8����E_^[���   ;��������]����������������������������������������������������������������������������U����   SVW��<����1   �������E���$��Y ��ٝ<���م<���_^[���   ;��e�����]����������������������������������U����   SVWQ��4����3   ������Y�M��E��E�X�M��E�Y�U��E��E�_^[��]� �����������������������U����   SVW��<����1   ������E� �E������Dz0�M�A�E������Dz�U�B�E������Dzǅ<���   �
ǅ<���    ��<���_^[��]�������������������������������������������U����   SVW��$����7   ������M�������̉�,���j h� ������$����M該���M�T����M�L������̉�8���j h� �̳����$����M�t���_^[���   ;�谶����]���������������������������������������������U��j�h~�d�    P��<  SVW�������O   ������XD3ŉE�P�E�d�    j h�.�M��/����E�    �EЫ� j h�.�����������E�j h�.������������E�j ������P������Qh~�j �U�R�E�P�z�����������������E��������#����E� ������������������t!ǅ����    �E������M�������������ǅ���   �E������M�����������R��P� �輨��XZ�M�d�    Y_^[�M�3�������H  ;��$�����]�   �����   �name �������������������������������������������������������������������������������������������������������U����   SVW��0����4   ������h�.jIhij�7�������8�����8��� t��8����n�����0����
ǅ0���    ��0���_^[���   ;��*�����]���������������������������������������U����   SVWQ��4����3   ������Y�M��M��i����E�� $/�E�_^[���   ;�蹳����]����������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P��������E�_^[���   ;��N�����]� ������������������������U����   SVWQ��4����3   ������Y�M��M�������E�� |/�E�_^[���   ;�������]����������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;�蕲����]������������������U����   SVWQ��4����3   ������Y�M��M������_^[���   ;��E�����]������������������U����   SVWQ��4����3   ������Y�M��M��P����E��t�E�P荥�����E�_^[���   ;��ޱ����]� ������������������������U��j�hʹd�    P��,  SVW�������  ������XD3ŉE�P�E�d�    �E�P�M�d�����������E�    �E�P�M��7����E�P�M�Q�M��Ǳ�����A  �M������P�M�迾���E���t���P�M�������E���t����������h�����P���P�M������E���P����������D�����h���P��h���+�D���Q��t����<�����,���P�M�n����E���,����}����� ����� ���P������Q�M�ǻ���������������������E��������@����� ���+�Q��,����ͨ���E�����������j h�/�������4����E�������P��,����A����E�������������t�����������&  ������P�M�߿�����u����E�j ������������E���P���P�� ���������E�	������Q�� ���R譱����������E��� ����/�������� �  ǅ����    ���������������������	��  ������P������Q�������E�
��t���P�����������������������������E�������R��P����?����E���P���P�������)����E�������Q��P���R������P������Q��������D����E��������S����E���P����D����E�
��t���������D��� ��   ������P�������X����������������������E�������R��t��������E�
����������������P�����������������������������E�����������P������R�������ۜ���������������������E�������谿��+�D���P��t����?����E��������)����E�
�����������E��������9�����E��������(��������  j h�/�������m����E�������P�����Q�������1����������������������E�������P��(���Q�2������������������������E�������P��t����=����E���(����^����E�������O����E��������@�����t���P��L���������E���P���Q��p���������E�������R��L���P��p���Q������R�ϝ�����������C����E���p��������E���L���������C�����tUj h�/�������7����E����ĉ�������P���Q������RP�������������M蹧���E��������e����E�������脠���E��������u������̉�������,���P�ø���������������������E����̉�������P���R薸���������������������E����̉�������t���R�i����������EP�E��c�����4�������������������E���,��������E���P��������E���t��������E� �M�裟�������E������M��H���R��P�h��T���XZ�M�d�    Y_^[�M�3��6�����8  ;�輪����]�   p�����   A�����   >�����   ;�����   7�����   4�t���   $�P���   �,���   �����   �����   ������   ��searchPath temp documentPath out bitmapFileName bitmapDirectory fn dat id bc ctr ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H�Q,�҃�;�蘧��_^[���   ;�舧����]� ����������������������������������U��j�h�d�    P��   SVW�������@  ������XD3ŉE�P�E�d�    �E�   �EP�MQ�U�R�������E��EP�M�������E��E�    j hL�M��٣���E��M��:�����u`ǅ ���    �E��M��$����E��M������E��M������E��M� ����E� �M������E������M,������ ����I  �M��8������E�y`ǅ���    �E��M�贾���E��M�訾���E��M�蜾���E��M萾���E� �M脾���E������M,�u����������  �EP��|��������E��M��������Ԫ�����E  ��d��������E��E,P��L���赲���E����̉�����EP蝲����������4���Q豠�����������E�	j h0������h����E�
�E�P������Y����E�j h �������?����E���L���P�������-����E�j h0�����������E��E�P������Q������R��$���P��������������������������E�������R��t���P�й�����E���$����$������̉�<�����t���P蠱���������n�������������������h������̉�H����E�P�l����������:�������������������\������̉�T���������P�5�����������������������������P���������P��P���Q耦������D�����D����u��P���P�
�������P���P�B�����ǅ8���    ǅ,���    ǅ ���    �M�������M�������������������������n'  t������o'  t������p'  t�"ǅ8���   �ǅ,���   �
ǅ ���   ǅ���    ǅ����    j j ��h���P�ɟ���������������� �Q  j j ��\���P裟���������������� �  ������P������Q�F�������t���P������Q�0�����������;�������   |������;�������   ��8��� u~��,��� uu��D��������E����̉�`���j ��\���P�[�����������D��������j j j�j���D���蝶����tǅ ���   �
ǅ ���    �E���D����A�����8��� t
ǅ���   �� ��� t
ǅ���   ������P�������
ǅ����   ������P�˭�����;j j ��\���P�R�������8�����8��� ~ǅ���   ��8���P莭��������� t!��j ��h���P��\���Q�T�;��[����(������ t��j ��\���P��h���Q�T�;��1�����P���P蔛������\���P腛�����E���t����s����E��������d����E��������U����E��������F����E�
������7����E�	������(����E���4��������E���L����
����E���d��������ǅl���   �E���|��������E��M��ָ���E��M��ʸ���E��M�辸���E��M貸���E� �M覸���E������M,藸����l���R��P�8�脓��XZ�M�d�    Y_^[�M�3��f�����  ;�������]�   @�����   ������   ������   ��|���   ��d���   ��L���   ��4���   �����   �����   ������   �����(  v�����   h�����   ^�t���   O�\���   D�P���   <�����0   7�t���0   2�D���(   $�confirmdialog sBuf dBuf destDir bitmapFile destFileString backSlash destDirString fileinfo space sourceFile slash wrlFileName destPath progressText path url fileName bitmapFileString ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hx�d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M�M�襵���E�    �E�� 0�M���ɣ���E������E�M�d�    Y_^[���   ;��f�����]���������������������������������������������������U��j�h��d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M��E�    �M���K����E������M��0����M�d�    Y_^[���   ;�貚����]�����������������������������������������������U����   SVWQ��4����3   ������Y�M��M�膾���E��t�E�P�ݍ�����E�_^[���   ;��.�����]� ������������������������U��j�h��d�    P��  SVW�������E   ������XD3�P�E�d�    ǅ����    �E�   j �M������P�m������������������E�j j �M������P�E�P�M������E�   �E�Ph`b艸�����E�`b�E������   �E������   �E���� ��   �E����'��   �E����"��   �E����\t�E����{tt�E����}ti�E����,t^�E����.tS�E����[tH�E����]t=�E����.t2�E����#t'�E����}�}� t�E����0|�E����9�E�� _�E�    �E����E������E쉅����������Q�u�����j h`b�M�J������������������E� �M蠰���ER��P�$�萋��XZ�M�d�    Y_^[��   ;�������]Ë�   ,�����   8�_$ArrayPad ���������������������������������������������������������������������������������������������������������������������������������������������U��j�h_�d�    P��  SVW�������D   ������XD3ŉE�P�E�d�    ǅ����    �E�   �E�    j �M�B����E܋�h@0�B��P�M܃�Q��c�B��H  �у�;�蹖���E�}� u*j �M�������������������E� �M������E�jj�E܃�P�M�Q�M�����E܋E�P�M�謡���E��E�P�Đ�����E�P�M荟�����������������E��M������E� �M莮���ER��P�@�~���XZ�M�d�    Y_^[�M�3��`�����  ;�������]Ë�   H����   j����    `StringSTD charline �������������������������������������������������������������������������������������������������������������U��j�h��d�    P���   SVW�������?   ������XD3�P�E�d�    �E�    �E�    j �M�?����E���h@0� B��P�M���Q��c�B��H  �у�;�趔���E�}� u!ǅ����    �E������M�����������6j�E���P�M�Q�M������E��E쉅����E������M�ˬ�������R��P��踇��XZ�M�d�    Y_^[��  ;��*�����]Ë�   ����   _$ArrayPad �������������������������������������������������������������������������������������U��j�h�d�    P��  SVWQ�������A   ������Y�XD3�P�E�d�    �M�M��V����E�    �M��@�D����E��M���   耛���E��M���   �n����E������M쉁�   j �M蚞���M쉁�   ������P�M�����������������������E�������R�M���   �����E��������1��������P�M蒁���������������������E�������R�M���   �ǭ���E�����������E�M���   �E�ǀ�       �E�ǀ�      �E������E�M�d�    Y_^[��  ;��.�����]� ��������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��c���_^[���   ;�腑����]������������������U��j�h�d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M��E�   �E��   P豏�����E��   P譇�����E��M���   �b����E��M���   �P����E� �M��@託���E������M�虗���M�d�    Y_^[���   ;�訐����]�����������������������������������������������������U����   SVWQ��4����3   ������Y�M��E����   _^[��]��������������U����   SVWQ��4����3   ������Y�M��E����   _^[��]��������������U����   SVWQ��4����3   ������Y�M��E����   ���U����   _^[��]������������������U����   SVWQ��4����3   ������Y�M��E����   ���U����   _^[��]������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �E��   P�M������,�������,����E_^[���   ;��������]� ��������������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �E��   P�M蔛����,�������,����E_^[���   ;��p�����]� ��������������������������U����   SVWQ��4����3   ������Y�M��E�ǀ�       _^[��]��������������������������U����   SVWQ��4����3   ������Y�M��E����   _^[��]��������������U��j�h��d�    P��D  SVWQ�������Q   ������Y�XD3�P�E�d�    �M��E�    �E싈�   �M��}� u$ǅ����    �E������M軥���������Z  �E�    j�M脄���Eȋ�h@0�$B��P�Mȃ�Q��c�B��H  �у�;�������Eԃ}� u$ǅ����    �E������M�H�����������   j�Eȃ�P�M�Q�M�6����EȋE샸�    t8�E�    �	�E����E��E�M�;��   }j �M�貛��j �M�訛������E�ǀ�      �E�    �	�E����E��E�;E�}9�E�E��Q�M��k�����u!ǅ����    �E������M苤���������-붍E�P�x�����ǅ����   �E������M�\���������R��P�l�I��XZ�M�d�    Y_^[��P  ;�軋����]� �   t����   �����   �_$ArrayPad charline ������������������������������������������������������������������������������������������������������������������������������������������������U��j�h�d�    P���   SVWQ������9   ������Y�XD3�P�E�d�    �M��E�   �M���ڒ���E��M��(�˒���E��E�E��M��u���M�A�M�蘌���M�A�M�踤���M�A�M��=����M�A�M蔓���M�A�EP�M���m����E�M��EP�M��(�V����E� �M�z����E������M�k����E�R��P�\�[}��XZ�M�d�    Y_^[���   ;��͉����]�$ �I    d����   p_$ArrayPad �������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�j h�  �M���s��_^[���   ;�������]���������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HH���  �҃�;�襈��_^[���   ;�蕈����]� �������������������������������U����   SVWQ��4����3   ������Y�M�h�  �M��t��_^[���   ;��0�����]�����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH���   �у�;��ȇ��_^[���   ;�踇����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�j h�  �M��
r��_^[���   ;��N�����]���������������������������U����   SVWQ��4����3   ������Y�M�h�  �M���r��_^[���   ;��������]�����������������������������U��j�hV�d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M��E�   �E�P襛�����E� �M��(�۞���E������M���ɞ���M�d�    Y_^[���   ;��?�����]��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �E���P�M�V�����,�������,����E_^[���   ;��2�����]� ����������������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �E���(P�M�֐����,�������,����E_^[���   ;�貃����]� ����������������������������U��j�h��d�    P���   SVWQ������6   ������Y�XD3�P�E�d�    �M��E�    �EP�M��(�w����E������M蘛��R��P�,�v��XZ�M�d�    Y_^[���   ;��������]� �I    4����   @_$ArrayPad �����������������������������������������������������U����   SVWQ������9   ������Y�M���#����̌��P��/�������P�M������E�_^[���   ;��J�����]�����������������������U��j�hӹd�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M��E�   �M�� �%����E� �M���߈���E������M��}���M�d�    Y_^[���   ;�裁����]������������������������������������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �EP�M����mu����,�������,����E_^[���   ;�������]� ����������������������������U����   SVWQ������;   ������Y�M�ǅ,���    ���ĉ� ���P�M��`���������MQ�UR�M��|����������,�������,����E_^[���   ;��q�����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M��M������j�M���i��_^[���   ;�������]���������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �EP�MQ�M��lk����,�������,����E_^[���   ;������]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�M�膢���������_^[���   ;������]� ���������������������������������U����   SVWQ��4����3   ������Y�M��M�袍��_^[���   ;��~����]������������������U��j�h�d�    P���   SVWQ������6   ������Y�XD3�P�E�d�    �M�EP�M���|���E�    �EP�M���|k���E��EP��#����ƚ����#���Q�M�� 資���E��E���0�X<j�M���g���E������E�M�d�    Y_^[���   ;���}����]� ������������������������������������������������������������������U��j�h��d�    P��8  SVWQ�������N   ������Y�XD3�P�E�d�    �M�ǅ ���    �EP�M�������E��M�袀���E�   �E�P�M�� �{��P������Q�M�訕���������������������E�������P�M��(n���E��������}����M��j����E�P�M���Q�M�� �z�����"���Ѕ��  �EP�M��;���P�'�����P�M���H����ȅ���   �M�����P�������P�EP�M�������ȅ�tB������R�M������������������������E��� ������� ����������������	�Ẻ�����������������������R�M袄���� ������� ����E�   �� �����t�� �����������h|���E� �M��\|���E�/������EP�M��C����� ������� ����E� �M��+|���ER��P����n��XZ�M�d�    Y_^[��D  ;��H{����]� ��   �����   �_Where ���������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h�d�    P���   SVWQ������:   ������Y�XD3�P�E�d�    �M썅���P�M����������������������E�    �����R�E��P�M�� �����E�����������z���E���M�A4�E�M�H8�M�d�    Y_^[���   ;��y����]� �����������������������������������������������������U��j�h��d�    P��  SVWQ��������   ������Y�XD3�P�E�d�    �M�ǅ����    �E�   �EP輋����P�M������E��E���P�M�� �
w��P�M�Q�M�藑���E��E�P�M�� ��v��P������Q�M��t����������������������E�������P�M��${���������E��������My�����������c  �M��n�����!���P������P�EP� �����P�M���!����ȅ�t�!  3�u1�EP�؊����P�M��ڟ��P�Ɗ����P�M�������ȅ�t�M�豚����   ��   �����P�M�訊���������������������E�������R�M�Hz��������E�������qx���������t=���̉�,����EP�dk����������8���Q�M���||����������8����)x��ƅO��� ��O���P�M�Q�M�������������������E��M���w���E� �M��w���E�o  �5�����d���P�M��ɉ���������������������E�������R�M�iy����[����E���d����w����[�����t\���̉�x����EP�j���������������������E��U��R���̉������E�P�Tj���������M���E��ff���d�EP���̉������U�R�%j��������������P�M���m���������������������E�������R�M�hg���E���������v���	�E����E��E�P�M�� � t��P������Q�M�芎���������������������E�������P�M������������E��������cv����������t'�EP�M�Q�M�� �s������f���}� u��l����M��~���M�ݝ�����k��ܝ��������AuY�M�� �{g����E��M��L����E��E�    �	�E����E��}�}�E�;E�s
�E����E��ߋE�P�M���^���M���|��ƅ����������P�MQ�M�u������������������E��M��u���E� �M�tu���ER��P��"�h��XZ�M�d�    Y_^[��$  ;��t����]� �I    �"����   �"_Plist ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U��j�h�d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M��E�    �M���`���E������M��s���M�d�    Y_^[���   ;��%r����]����������������������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �E�P�M��QR�M�˄����,�������,����E_^[���   ;��q����]� ����������������������������������������U����   SVWQ������9   ������Y�M�j �E�P�M��Ő���E��HQ�ve������U��E��HQ�be�����U��J��E��HQ�ݑ�����U��J��E��@    ��E�E��E��M�;Ht3�E�P�e������M�E�P�M����Ȇ��j�E�P�M��������_^[���   ;��p����]����������������������������������������������������������U��j�h�d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M��E�    �M��6����E������M��2����M�d�    Y_^[���   ;���o����]����������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��Tk���E��M�P3�;Q��_^[���   ;��po����]� ��������������������������U����   SVWQ��4����3   ������Y�M��EP�M������E�_^[���   ;��o����]� ������������������������U����   SVWQ��4����3   ������Y�M��EP�M��b���E�_^[���   ;��n����]� ������������������������U����   SVWQ��4����3   ������Y�M��EP�M�肉���E��M�Q�P�E�_^[���   ;��Bn����]� ����������������������������U����   SVWQ��4����3   ������Y�M��M��s���_^[���   ;���m����]������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��m����]������������������U����   SVWQ��4����3   ������Y�M��EP�M���|���E��M�Q�P�E�_^[���   ;��2m����]� ����������������������������U����   SVWQ��4����3   ������Y�M��EP�M��"����E�_^[���   ;���l����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��^��_^[���   ;��ul����]������������������U����   SVWQ��4����3   ������Y�M��EP�M��=����E�_^[���   ;��l����]� ������������������������U����   SVWQ��4����3   ������Y�M��EP�M��&]���E�_^[���   ;��k����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��;n��_^[���   ;��ek����]������������������U����   SVWQ��4����3   ������Y�M��EP�M��>l���E�_^[���   ;��k����]� ������������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �EP�M�rs����,�������,����E_^[���   ;��j����]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��@8_^[��]�����������������U����   SVWQ������:   ������Y�M��M��gS����,���ǅ0���    ߭,����M�ݝ$������������ǅ ���    ߭���ܽ$���ٝ���م���_^[���   ;��i����]��������������������������������������U����   SVWQ��4����3   ������Y�M��E��@<_^[��]�����������������U����   SVWQ��(����6   ������Y�M��EP�M����[����M�#A4�E�E��H8;M�w�E��H4����U�+щU�E�_^[���   ;���h����]� ������������������������������U��j�hi�d�    P��H  SVWQ�������R   ������Y�XD3�P�E�d�    �M�M���k���E�    j �M�� �Yf��P������P�M������������������������E�������R������P�M����^���������������������E�������R�M��4Y�����]j���������E��������h���E� �������wh����������t\���̉������E�P�_p���������������������E��M��,���P�� ���R�E� �M��U���������� ����c[��������E������M��h��R��P�0�Z��XZ�M�d�    Y_^[��T  ;��!g����]Ð   0����   0_First �����������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��t���E��U��J�E�_^[���   ;��Gf����]� ���������������������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M��XV��_^[���   ;��e����]� �����������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��@����0   ������E��_^[��]����������������������U��j�h��d�    P���   SVWQ������6   ������Y�XD3�P�E�d�    �M�Q�̉� ����EP�e���M���i���E�    �M��݀���M�A�E��@    �E������E�M�d�    Y_^[���   ;��`d����]� ������������������������������������������U��j�h��d�    P���   SVWQ�������>   ������Y�XD3�P�E�d�    �M�ǅ ���    �E�   �EP���̉�����UR�W���� ����M��|���M�Z�����̉����P�dW���� ����EP�M��i���������� ������� ����E� �M�q���E�M�d�    Y_^[��  ;��Mc����]� �����������������������������������������������������������������������U��j�hb�d�    P��  SVWQ�������C   ������Y�XD3�P�E�d�    �M�ǅ���    �E�   �E;E�u�E�M;Huh  h�"h�"�{����j ������P�M袂���������������������E��������G{���E��E��������^p���E�P�M�Q�M�赁���E�M�;H��   �E�P�ZV�������M�Q�ނ�����R�AV�������E�P�Â�������M�Q�#V�����R誂�������E�P�M����w��j�E�P�M����s���E�H���U�J���̉�����EP�QU���������MQ�M���f���������������������E� �M�wo���E�M�d�    Y_^[��  ;��:a����]� ��������������������������������������������������������������������������������������������������������������������U��j�hٽd�    P��8  SVWQ�������N   ������Y�XD3�P�E�d�    �M��E�   ������P�M�T���������������������E�������R�M蘃���������E���������`����������thw  h�"h�0�Fy������   �EP�M���S���E��M��L����E�;Eu.�EP�M�Qb���ȅ���   �E�P�M�:b���ȅ���   j j���̉������E�P�gS���������������������E����̉� ����UR�=S���������������������E��MQ���̉�����UR�S���������E��M�� l���E��M��Jm���E� �M�>m���E������M�/m��R��P�D8�rR��XZ�M�d�    Y_^[��D  ;���^����]� ��   L8����   X8_Last ����������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M���b���E��HQ�LR����P�M����#����E��HQ��~����P�M�������j�E��HQ�M�����o���E��@    _^[���   ;��]����]����������������������������������������������U����   SVWQ������9   ������Y�M�j�M��([���E�E��E��8 tJ�E���U��A;Bt�} t�E���Q;Ut�E�����M���E���    �E���U��A�뮍M�超��R��P�T:�UP��XZ_^[���   ;���\����]�    \:����   h:_Lock ������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��"k��_^[���   ;��5\����]������������������U����   SVWQ��4����3   ������Y�M��EP�O����_^[���   ;���[����]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�K����_^[���   ;��[����]� ���������������������������U��j�h�d�    P���   SVWQ������6   ������Y�XD3�P�E�d�    �M�Q�̉� ����EP�a���M���f���E�    j �M��K���E������E�M�d�    Y_^[���   ;���Z����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��M�����G��_^[���   ;��bZ����]�������������������������������U����   SVWQ��4����3   ������Y�M��M��[s��;EwZh  hP6h6�3s����3�u!h�$j h  hP6j��K������u�j h  hP6h81h�#�_�����M���r��9ErC3�u!h1j h  hP6j�xK������u�j h  hP6h81h�#�^_����3�u��Ek��M�A_^[���   ;��FY����]� ����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M���M��_^[���   ;��X����]� �����������������������U����   SVWQ��4����3   ������Y�M��E��x tE�M���X���E��HQ�U��BP�M��Q���E��M��@+A��   ��P�U��BP�M�����\���E��@    �M��A    �U��B    _^[���   ;��X����]����������������������������������������������U����   SVWQ��4����3   ������Y�M��M��f��_^[���   ;��W����]������������������U����   SVWQ��4����3   ������Y�M��M��Q���E�_^[���   ;��BW����]�������������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M��~���E�_^[���   ;���V����]� ��������������������U����   SVWQ��4����3   ������Y�M��M��7U��_^[���   ;��V����]������������������U����   SVWQ��4����3   ������Y�M��M�袀���E�_^[���   ;��2V����]�������������������������������U����   SVWQ��4����3   ������Y�M��M��DL���E�_^[���   ;���U����]�������������������������������U����   SVWQ��4����3   ������Y�M��E��8 t�E��M�;tch<  h�"h�)�n�����   ��tC3�u!h@)j h=  h�"j�(G������u�j h=  h�"h�6h$(�[����_^[���   ;��U����]� ������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��\]���E��M��P�E�_^[���   ;��T����]� �����������������������������U����   SVWQ��4����3   ������Y�M��M����h��_^[���   ;��"T����]�������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVWQ������>   ������Y�M��EP�g����%����E�h� �E�P�a��������������������M܋�����U��E�i��A  �M�i�  +��E�y�E�����E��E�R��P�D�F��XZ_^[���   ;��S����]�    D����   (D_Qrem ������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�RX����_^[���   ;��mR����]� �����������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �E�P�M��QR�VF����� P�M�e����,�������,����E_^[���   ;���Q����]� �����������������������������U��j�hg�d�    P���   SVWQ������6   ������Y�XD3�P�E�d�    �M�ǅ ���    �E�   �E�P�MQ�M�hd���� ������� ����E� �M�a_���E�M�d�    Y_^[���   ;��$Q����]� ����������������������������������������������U��j�h��d�    P���   SVWQ������9   ������Y�XD3�P�E�d�    �M��E�    �E;E�th�  h�"h�#��i�����M�vi���E��EP�M�Q�Eq�����R�E�P�M��{L���E�j�M���n���E�P�q�����Mԉ�E�P�q�����Q�oD�����Uԉ�E������M�4^���M�d�    Y_^[���   ;���O����]� ��������������������������������������������������������������������U��j�h�d�    P��d  SVWQ�������Y   ������Y�XD3�P�E�d�    �M��E�   �E;E�thi  h�"h�0�h�����E��P�M��Q��R�����Ѕ���  �E4����   �E�;Et}�EP�M���B���E��E$P�M��mQ���ȅ�tNj ������P�M��o���������������������E��������BP�MQ�M��9n���E���������\����E��M��\���E�;Et�E0P�M��m���E�H+M0�U�J�M$�ag�����M�Wg��P�0o����� P�B�����0�M�9g�����M$�/g��P�o����� P�kB�����0�M�g�����M�g��P��n����� P�CB�����0�M��f��P��n����� �E̍M$��f��P�n�������M��f��P�n�������M�f��P�n�������M$�f��P�qn�������M�f��P�\n�����M̉��   ���̉������E$P�,A���������������������E����̉������UR�A���������������������E����̉������UR��@���������E��M���6�����̉������E$P�@���������������������E����̉������UR�@��������������P�E��M�XH���������������LM���E��M�Z���E� �M�Z���E������M$�Z��R��P��J��?��XZ�M�d�    Y_^[��p  ;��EL����]�0 �I    �J����   �J_Next ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h`�d�    PQ���   SVWQ������:   ������Y�XD3�P�E�d�    �e��M�j�M���I���E��E�    �E�    �E�P�?����������M�Q�����R�M���Z���EЃ��EЋE�P�gk����������M�Q�����R�M���|Z���E�}� ~�E�P�>����P�M���|l��j�E�P�M���v\��j j �xo���E�������L��E������E�R��P�0M�=��XZ�M�d�    Y_^[���   ;���I����]Ë�   8M����   DM_Pnode �����������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M�Q�̉�,����EP�I���M��'s���EP�M����yI���E�_^[���   ;��I����]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�B����_^[���   ;��H����]� ���������������������������U����   SVWQ��4����3   ������Y�M��E��M��@+A��   ��_^[��]�������������������U��j�hĿd�    P��t  SVWQ�������]   ������Y�XD3�P�E�d�    �M�EP�M��P���E�    ������P�M��SN���������������������E����̉�����������R�Z���������������������E�������Q�M���A���������������������E����̉�����������P��Y��������������Q�E��M��}Y����������������R���E���������R���E� ��������R���E�P�MQ�����R�M��TA���������������������E����̉�����������R�AY���������M��:4���E� ������R���E������M��YG��R��P��P�:��XZ�M�d�    Y_^[�Ā  ;��yF����]� �I    �P����   �P_Tmp ���������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@    �M��A    �U��B    �} u2��K�G�M��7��;Es�:���3�EP�M����K<���M��A�E��M��Q�P�Ek��M�A�U��B�_^[���   ;��*E����]� ����������������������������������������������������U����   SVWQ��4����3   ������Y�M��E���P�MQ�UR�d����_^[���   ;��D����]� ��������������������������������U����   SVWQ��(����6   ������Y�M�Q�̉�,����EP��J���M���:���EP�M����J���E�_^[���   ;��!D����]� ���������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVWQ��4����3   ������Y�M��EP�-7����_^[���   ;��C����]� ���������������������������U����   SVWQ��$����7   ������Y�M��E�UUU�}� v�E쉅$����
ǅ$���   ��$���_^[��]�������������������������������U����   SVWQ��4����3   ������Y�M��M��+-���E��@    �E�_^[���   ;��B����]���������������������U��j�h�d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M�M��,���E�    �E�M�H�EP�M��A���E������E�M�d�    Y_^[���   ;��B����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 t�E��x t�E���U��B;Auch�   h�"hX%�Z�����   ��tC3�u!h�$j h�   h�"j�;3������u�j h�   h�"h89h�#�!G�����E��HQ��]����_^[���   ;��
A����]�������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 t�E��x t�E���U��B;Auch�   h�"h�&�Y�����   ��tC3�u!h�$j h�   h�"j�;2������u�j h�   h�"h�;h�#�!F�����E��HQ�`4�����U�� �B�E�_^[���   ;���?����]������������������������������������������������������������U��j�hW�d�    P���   SVWQ������;   ������Y�XD3�P�E�d�    �M�ǅ���    �E�P�M��.3���E�   �M��i���E�P�M�3���������������E� �M��QM���ER��P�$X�2��XZ�M�d�    Y_^[���   ;��?����]� �   ,X����   8X_Tmp �������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 t0�E��x t'�E��HQ�5_�����U�� �B�M���E��H;Juch  h�"h�'�hW�����   ��tC3�u!h�$j h  h�"j��/������u�j h  h�"h�=h�#��C�����E�_^[���   ;���=����]������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��M��|J��_^[���   ;��=����]������������������U����   SVWQ��4����3   ������Y�M��EP�M��n;���E��M�Q�P�E�_^[���   ;��<����]� ����������������������������U����   SVWQ��4����3   ������Y�M��M��m>��_^[���   ;��U<����]������������������U����   SVWQ��4����3   ������Y�M��M��tK���E�_^[���   ;��<����]�������������������������������U����   SVWQ��4����3   ������Y�M��EP�M���Z���E�_^[���   ;��;����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��<��_^[���   ;��E;����]������������������U����   SVWQ��4����3   ������Y�M��M��}T���E�_^[���   ;���:����]�������������������������������U����   SVWQ��4����3   ������Y�M��EP�M���+���E�_^[���   ;��:����]� ������������������������U����   SVWQ��4����3   ������Y�M��M���Q��_^[���   ;��5:����]������������������U����   SVW��@����0   ������E��_^[��]����������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U��j�h�d�    P��L  SVWQ�������S   ������Y�XD3�P�E�d�    �M�ǅ ���    �E�   ������P�M��0���������������������E��� ������� ���������P�M�_\���ȅ�tY������R�M��--���������������������E�   �� ������� ���������R�M�\������tǅ����   �
ǅ����    �������������E�   �� �����t�� �����������$9���E�   �� �����t�� ����������� 9����������tH�M���<���EP�M��f,���� ������� ����E��M�1F���E� �M�%F���E��   ��   �EP�M�c:���ȅ�t_���̉������EP�+���������� ���Q�M��<���������������������E�������P�M�\_���E��� ����=8��뎃��̉�����EP�9+���������MQ�M���<���������� ������� ����E��M�_E���E� �M�SE���E��E��M�BE���E� �M�6E���M�d�    Y_^[��X  ;���6����]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h`�d�    PQ���   SVWQ������:   ������Y�XD3�P�E�d�    �e��M�j�M����4���E��E�    �E�    �E�P�*����������MQ�����R�M���E���EЃ��EЋE�P�wV����������MQ�����R�M���E���EЃ��EЋE�P�,R����������MQ�����R�M���A2���c�}�~�E�P�V����P�M���[W���}� ~�E�P�f)����P�M���=W��j�E�P�M���7G��j j �9Z���E������:b��E������E܋M�d�    Y_^[���   ;���4����]� ��������������������������������������������������������������������������������������������������U��j�h��d�    P��(  SVWQ�������J   ������Y�XD3�P�E�d�    �M�M���"���M�+A;EsLh�)������E?���E�    �����P�������`G��h��������Q�Y���E�����������2���E�HM�U�J�M�d�    Y_^[��4  ;��3����]� ���������������������������������������������������������������U����   SVWQ��(����6   ������Y�M�Q�̉�,����EP�p3���M��N���EP�M����A(���E�_^[���   ;���2����]� ���������������������������U����   SVWQ��4����3   ������Y�M�j �EP�X;����_^[���   ;��2����]� �������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�F����_^[���   ;��-2����]� �����������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �E�P�M��QR�M�\-����,�������,����E_^[���   ;��1����]� ����������������������������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �E�P�M��QR�M��,����,�������,����E_^[���   ;��1����]� ����������������������������������������U��j�h��d�    P���   SVWQ������7   ������Y�XD3�P�E�d�    �M��E�    �EP�MQ���̉� ����UR��B��������M��8���E������M��=���M�d�    Y_^[���   ;��S0����]� ���������������������������������������������U��j�h?�d�    P��,  SVWQ�������K   ������Y�XD3�P�E�d�    �M�ǅ����    �E�   ���̉������EP�)B���������M�Q�M��?���������E����̉������EP��A���������M�Q�M���>���������E��E�P�M��k4���ȅ���   �E�P�M��x���ȅ�u�E�;E�u�E�M�;Hr�E�H;M�sh  hP6h @�HH�����E�P�M�QR�E�P�UL�����E��E�HQ�U�R�M��:D���E�HQ�U�R�M��%(���E�M��H�E�P�M�Q�M�A*�����������������E��M��f:���E��M��Z:���E��M��;���E� �M��;���ER��P��h��!��XZ�M�d�    Y_^[��8  ;��G.����]� �   �h����   i����    i_Last _First �����������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P��  SVW�������G   ������XD3�P�E�d�    hx@������8���E�    �����P�������@��h��������Q�XR���E������������+���M�d�    Y_^[��(  ;���,����]���������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��:���E�_^[���   ;��r,����]� ����������������������������U����   SVWQ��4����3   ������Y�M�j �EP�)����_^[���   ;��,����]� �������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ������_^[���   ;��+����]� �����������������������U����   SVWQ��4����3   ������Y�M��M����H��_^[���   ;��R+����]�������������������������������U����   SVWQ��(����6   ������Y�M�Q�̉�,����EP�P+���M��T���EP�M����+���E�_^[���   ;���*����]� ���������������������������U��j�h��d�    P���   SVWQ������6   ������Y�XD3�P�E�d�    �M�ǅ ���    �E�   �E�P�MQ�M��%���� ������� ����E� �M�7���E�M�d�    Y_^[���   ;��*����]� ����������������������������������������������U��j�h8�d�    PQ��4  SVWQ�������M   ������Y�XD3�P�E�d�    �e��M��E�    �E;E�u�E�M;Hr�E�H;Msh�  hP6h�@�B�����M��f#���E܃} u�  �M��B�����M��b��+�;Es
�S���  �M��cB��E9E���  �u���M��0��+�;E�sǅ����    ��E���E܉������������M܋M��B��E9E�s�M��B��E�E܋E�P�M������EЋE�M+H����   ���E��E�    �E��EP�MQ�U�k�U�R�M���A���E����E��E�P�MQ�U�BP�M��;2���E����E��E�Ek�E�P�M�QR�EP�M��2���o�}�~�E�k�E�P�M�Q�M��_!���}� ~$�Ek��M�k�M��Q�U�k�U�R�M��5!���E�P�M�Q�M���,��j j �M���E�    �ro��E�    �M���@��E�E�E�x t=�E�HQ�U�BP�M��� ���E�M�@+A��   ��P�U�BP�M���,���M��'���E�k�EЋM�A�Ek�EЋM�A�E�MЉH�  �E�@+E��   ��;E��   �EP�M��/���E��Ek�EP�M�QR�EP�M���0���E��E�P�M�A+E��   ���U+�R�E�HQ�M��@���5�Ek��M�AP�Uk�UR�M�����j j ��K���E�   ��p��E�   �Ek��M�A�U�B�E�HQ�UR�M��;���E�P�Mk��U�B+�P�MQ�b2�����E� �M���&���   �EP�M���.���E��E�H�M��E�HQ�U�R�Ek��M�+�Q�M���/���U�B�E�HQ�UR�M��&;���E�P�Mk��U�+�R�EP�*�����E�P�Mk�MQ�UR��1�����E� �M��?&���E������M��2��R��P��q����XZ�M�d�    Y_^[��D  ;��P%����]� ��   �q����   �q����   �q_Tmp _Tmp ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ������9   ������Y�M�j�M��!���E��E��E��8 tA�E���Q;Ur�E���U;Qs�E�����M���E���    �E���U��A�뷍M��L��R��P��s���XZ_^[���   ;��;#����]� �   �s����    t_Lock ����������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M������E�_^[���   ;��"����]� ��������������������U����   SVWQ��4����3   ������Y�M��EP�M��B���������_^[���   ;��7"����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��EP�M�����E��M�P;Q���_^[���   ;���!����]� ���������������������������U����   SVWQ��$����7   ������Y�M��E�����}� v�E쉅$����
ǅ$���   ��$���_^[��]�������������������������������U����   SVWQ��4����3   ������Y�M��M��)/���E�_^[���   ;��� ����]� ����������������������������U����   SVWQ��0����4   ������Y�M��E��x uǅ0���    ��M��U��A+B��   ����0�����0���_^[��]����������������������������������U����   SVWQ��4����3   ������Y�M��E���P�MQ�UR�EP�F�����Ek�E_^[���   ;�������]� �����������������������������������U��j�hx�d�    P���   SVWQ��(����3   ������Y�XD3�P�E�d�    �M�M���/���E�    �} tS�E�H;Mw�E�M;Hv=3�uh�Ej jFhP6j�5������u�j jFhP6h�@h$(�%����3�u��EP�M������E�M�H�E������E�M�d�    Y_^[���   ;�������]� ������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M�����E��M�P3�;Q��_^[���   ;��P����]� ��������������������������U����   SVWQ��4����3   ������Y�M��E��8 t�E��M�;tZh�   hP6h�K�7����3�u!h@)j h�   hP6j�������u�j h�   hP6h Gh$(�#����_^[���   ;������]� �����������������������������������������U����   SVWQ��4����3   ������Y�M��M�����E�_^[���   ;��"����]�������������������������������U����   SVWQ��4����3   ������Y�M��M��M6���E�_^[���   ;�������]�������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVW��@����0   ������j �M�8&��_^[���   ;��(����]���������������������U����   SVW��4����3   ������M�T���E��M�!��E�P�E�P��C����_^[���   ;������]����������������������������U����   SVW��4����3   �������E�ŝ��E;Et�E�i�� �M�3E��E���E�ًE�_^[��]���������������������������U����   SVW��@����0   ������EP�M���3Ʌ�����_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M��M����P�M�J!��P�E��HQj �M����_^[���   ;��z����]� ������������������������������������U����   SVWQ�� ����8   ������Y�M��} th�  h0*�EP�������E��H;Ms�=���E��H+M;Ms�E��H+M�M�E;Es�M��$����	�U��$�����$���P�MQ�M��f ��EP������E�}� t�E쉅$����1�M;Msǅ ���������U3�;U���� ����� �����$�����$���_^[���   ;��Q����]� ���������������������������������������������������������������������������U����   SVW��@����0   ������EP�MQ�UR�!����_^[���   ;������]���������������������������U����   SVW��@����0   ������_^[��]����������U��j�h��d�    P��  SVWQ�������G   ������Y�XD3�P�E�d�    �M��E�   �EP������Q�:����������R���̉�����E P����������������������E����̉�����UR����������������������E����̉� ����UR�j���������E��M��?���E��M�%���E� �M�%���E������M �%���M�d�    Y_^[��(  ;��P����]�$ ��������������������������������������������������������������������������U����   SVW��@����0   ������_^[��]������������U����   SVW��4����3   ������EP�MQ�7������;�����;���R�EP�MQ�UR�����_^[���   ;��p����]�����������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVW��,����5   ������} w	�E    �+���3��u��(sj ��0����X,��h<���0���P��:���Ek�(P�\����_^[���   ;������]��������������������������������������U����   SVW��$����7   ������E�E��E�Pj��*������,�����,��� t��,����U����,�����$����
ǅ$���    _^[���   ;�������]���������������������������������������U����   SVW������9   ������3���#����MQ�UR�5������/�����#���P��/���Q�UR�EP��;���Q������R�EP�MQ�����P�UR�����P��*����_^[���   ;��3����]������������������������������������������������U����   SVW��,����5   ������} w	�E    �+���3��u��sj ��0����H*��h<���0���P��8���Ek�P�L����_^[���   ;������]��������������������������������������U��j�h�d�    P���   SVW������:   ������XD3�P�E�d�    �E�E�E�Pj �(������ ����E�    �� ��� t�MQ�� ����1��������
ǅ���    �����������E������M�d�    Y_^[���   ;������]�������������������������������������������������������U����   SVW��@����0   ������_^[��]������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVWQ��4����3   ������Y�M��E���P�MQ�UR�EP�8����_^[���   ;������]� ����������������������������U����   SVW��@����0   ������EP�MQ�	����P�UR�	����P�����_^[���   ;��<����]�������������������������U����   SVW������9   ������3���#����MQ�+;������/�����#���R��/���P�MQ�UR��;���P�������Q�UR�EP������P�MQ������P������_^[���   ;������]����������������������������������������������������U����   SVW��(����6   ������3���/����MQ�UR�1������;�����/���P��;���Q�UR�EP�MQ�UR�w����_^[���   ;�������]�����������������������������������������U����   SVWQ��4����3   ������Y�M��M��/���E��t�E�P������E�_^[���   ;��^����]� ������������������������U����   SVWQ��4����3   ������Y�M��M������_^[���   ;������]�������������������������������U����   SVW��4����3   ������ER��P�|��!��XZ_^[��]ÍI    ������   ��_Cat ���������������������������U��j�hs�d�    PQ��D  SVWQ�������Q   ������Y�XD3�P�E�d�    �e��M��E�   h�  h�"���̉������E P�����������������������E����̉������UR����������E������� �EP�M�����E��E���M�8���E P�M�����������������t9�M�(��������������P���̉������UR�+���������M��/&����   ��M��7���EP�M�����ȅ�t]�EP�M��� ���E��M��z�����̉�����P�� ��������������P�M���������������������E��M������j j �2���E�   �g���E�   �E��M������E��M�����E� �M����E������M ���R��P�̊�����XZ�M�d�    Y_^[��T  ;��Z����]�(    Ԋ����   �����   �_Before _Next ������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��4����3   ������E�R��P�̋�����XZ_^[��]ÍI    ԋ����   ��_Cat ���������������������������U����   SVW��@����0   �������	�E���E�E;Et�EP�M������_^[���   ;���
����]������������������������������U����   SVW��4����3   �������E�P�MQ�G$����R��P�Č�����XZ_^[���   ;��`
����]�   ̌����   ،_Base_tag ������������������������������U����   SVW��4����3   ������ER��P�<��a���XZ_^[��]ÍI    D�����   P�_Cat ���������������������������U����   SVW������<   ������E+E��   ��k�E�E�3������3Ɉ�#��������R��#���P��/���Q�UR�����P�EP�MQ��)�����E�_^[���   ;��#	����]������������������������������������������������U����   SVW��(����6   ������3���/����MQ��2������;�����/���R��;���P�MQ�UR�EP�� ����P�MQ�� ����P�2����_^[���   ;��n����]�������������������������������������������U����   SVW��@����0   ������hU  h��EP�MQ�8&�����	�E���E�E;Et�EP�M�/�����_^[���   ;�������]������������������������������������U����   SVW��4����3   ������E�R��P��������XZ_^[��]ÍI    ������   ��_Cat ���������������������������U����   SVW��(����6   ������3���/����MQ�UR� (������;�����/���P��;���Q�UR�EP�MQ�UR�����_^[���   ;�������]����������������������������������������U��j�h��d�    PQ���   SVW��$����3   ������XD3�P�E�d�    �e��E�E��E�    ��E���E�M���M�} v�EP�MQ�M�,�����7�	�E���E�E�;Et�E�P�M������j j �9+���E������:���E������M�d�    Y_^[���   ;�������]��������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�r�����_^[���   ;��M����]� �����������������������U����   SVWQ��4����3   ������Y�M��EP�#����_^[���   ;�������]� ���������������������������U��j�h��d�    P���   SVW�������?   ������XD3�P�E�d�    �E�   �EP�����Q��&���������R�E$P�M Q���̉� ����UR������ ����� ����������E����̉�,����UR������������E��������$�E� �M�,���E������M����M�d�    Y_^[��  ;�������]����������������������������������������������������������������U����   SVW��@����0   ������E� _^[��]�����������������������U����   SVW��@����0   ������h�	  h��EP�MQ�X!������E���E�M���M�E;Et�EP�M�F����؋E_^[���   ;�������]����������������������������������������U����   SVW��@����0   ������EP�MQ�UR�EP�c����_^[���   ;��z����]�����������������������U����   SVW��4����3   ������EP��;���Q�r+�����R�EP�MQ�UR�EP�����_^[���   ;������]��������������������������������U����   SVW������<   ������E+E��   ��k��U+ЉU�3������3Ɉ�#��������R��#���P��/���Q�UR������P�EP�MQ�k*�����E�_^[���   ;��Q����]����������������������������������������������U��j�hD�d�    P���   SVW������:   ������XD3�P�E�d�    �E�E�E�Pj�X������ ����E�    �� ��� t�MQ�� ����e	��������
ǅ���    �����������E������M�d�    Y_^[���   ;��j ����]�������������������������������������������������������U����   SVW��@����0   ������j �M����_^[���   ;��������]���������������������U����   SVWQ��4����3   ������Y�M��M��i ���E��t�E�P�=������E�_^[���   ;�������]� ������������������������U��j�hx�d�    P���   SVW��4����0   ������XD3�P�E�d�    �E�    �M�C���E������M�4���M�d�    Y_^[���   ;��������]���������������������������������������U����   SVW��(����6   ������3���/����MQ�UR�������;�����/���P��;���Q�UR�EP�MQ������P�UR������P�
����_^[���   ;��J�����]���������������������������������������U����   SVW��4����3   ������ER��P�<��a���XZ_^[��]ÍI    D�����   P�_Cat ���������������������������U����   SVW��@����0   ������E;EtE�EP�MQ�UR��������EP�MQ�UR�������E;Es�EP�MQh4L�����_^[���   ;��5�����]����������������������������������U����   SVW��@����0   ������hr
  h��EP�MQ������E;Et �E���E�M���M�UR�M������؋E_^[���   ;�������]������������������������������������������U��j�h��d�    PQ���   SVW��$����3   ������XD3�P�E�d�    �e�j}hpL�EP�MQ�H����j~hpL�EP�T������E�E��E�    ��E���E�M���M�E;Et�EP�MQ�M�<"�����7�	�E���E�E�;Et�E�P�M�_�����j j �� ���E����������E������E�M�d�    Y_^[���   ;��l�����]�������������������������������������������������������������������������U����   SVW��@����0   ������} u�EP�MQh�*�!����_^[���   ;��������]��������������������U��j�h�d�    P��T  SVWQ�������U   ������Y�XD3�P�E�d�    �M�j h`M�������j����E�    ������P�M��*���E��������������j hHM�������0����E�   j hM�����������E�j ������P�M��Q������R������P�������������������������E�������R�����P�������������������������E�������Rj j j h�� �M��"���E�����������E������������E������������E���������������j�M������   �M�d�    Y_^[��`  ;��*�����]�������������������������������������������������������������������������������������������������������U��j�hH�d�    P���   SVWQ������6   ������Y�XD3�P�E�d�    �M��E�    �EP�M������E������M����R��P�������XZ�M�d�    Y_^[���   ;��-�����]� �I    �����   �_$ArrayPad �����������������������������������������������������U����   SVWQ��4����3   ������Y�M�j j hi'  �M��������u3���   _^[���   ;�������]����������������������������U���l  SVWQ�������[   ������Y�M�hl'  �������#���j j������P�M�����hm'  ������� ���h���h   �j jh���h   �hn'  ������P�M��H ��hq'  �����������j j������P�M��U���hv'  ����������h���h   �j jh���h   �hw'  ������P�M������hz'  �������e���j j ������P�M������h{'  �������B���j j ������P�M������hs'  ����������j j Q���$Q���$haerfQ��M�$Q���$Q���$Q�|M�$������P�M��) ��h}'  ����������j j�����P�M��\���h'  ���������j j Q���$Q���$haerfQ���$Q�xM�$Q�tM�$Q�pM�$�����P�M����ht'  ��(����P���j j��(���P�M�������   _^[��l  ;��2�����]�����������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��M��E��@    �E�_^[��]� �������������������������������U���l  SVWQ�������[   ������Y�M�hl'  �����������E���P������Q�M��	��hm'  ������������E���P������Q�M��I���hq'  �����������E��� P������Q�M�����hv'  �����������E���$P������Q�M������hz'  �������k����E���(P������Q�M��w��h{'  �������E����E���,P������Q�M��Q��hs'  �����������E���0P������Q�M�����h}'  �����������E���4P�����Q�M����h'  �����������E���8P�����Q�M����ht'  ��(��������E���<P��(���Q�M����3�_^[��l  ;�������]����������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@ _^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@$_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@(_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@,_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@0_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@4_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@8_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@<_^[��]�����������������U��j�h��d�    P���  SVW�� �����   ������XD3ŉE�P�E�d�    �} ��  �M��T����E�E�E�E܋M�}�����̉�@���P������8����E�P�2�������4����E�    �E�    �E�P��h���������E�������P�M��@�����8�����8�����4����E���4���R���̉�X�����h���P������0�����d���Q�(������,�����,�����(����E���(���P������Q�M��@�Q�����$�����$����� ����E��� ���������O����E�������������E���d��������E�������������O�������   j h�-������������E��E�P������Q�������8�����8�����4����E���4���P������Q�U�R������P�������0�����0�����,����E���,���R������P�s������(�����(�����$����E���$���R��h����~���E�����������E�����������E�����������E��������r���E����E�������h���P�M��%�����̉�����E�P�������8����� ���Q�`������4�����4�����0����E�	��0���P��H���Q�M��@�������H��������E��� ����f������̉�`���j h �[�����8����M����ǅ\���    �M�
�����P����M� �����D����M�5����������t
ǅP���    �M������	����t
ǅD���    ��P��� u��D��� u
ǅ\���   ��P��� u��D���u�} t
ǅ\���   ��P���u�} t��D��� u
ǅ\���   ��P���u�} t��D���u�} t
ǅ\���   ��\��� ��   �M�������tm�} u�EP�������E���̉�l����E�P�'�����8����MQ�UR����������̉�x����E�P�������8����MQ�UR�EP�������E�   �E�   ��E�    �E�    �EP�M�Q�U�R�M����P�EP�MQ��������M�����E�E� ��h��������E������M������ ���R��P�������XZ�M�d�    Y_^[�M�3��������  ;��:�����]Ë�   ������0   4�����   &�h���   �knotennametmp knotennameC4D mg �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�ha�d�    P��  SVW��T����h  ������XD3�P�E�d�    �E�    ���]����]��M�>�����
���]ԍE�P�M�������3����E�P�M��������S����E�P�M�Q�U�R��������M�������]�j hhN������������E�j h  �����������E����􉥔���������P�MQ������R������P�������������������������E�������RV�i������������M�����E������������E������������E� �������������̉�����j h`N�	����������M�����M�����E�    �	�E����E��E��E��X.������A��   �E��E��u����u��]�j h\N�� ��������E����������� ���Pj0j j�j�Q�E��$�����Q�.������������������������E�������PV�Y������������M������E�����������E� �� ��������E���   ����u+�}� t%���̉�0���j h ������������M����������M�A�����̉�<���j hXN������������M�i������̉�H���j hHN�����������M�D����M�D����E��X.ٽ����������   ������٭����߽����٭����������3ɺ   �������Q��������T�����T����E��E��X.ٽ����������   ������٭����߽����٭����������3ɺ   �������Q�������`�����`�����t����E��X.ٽ����������   ������٭����߽����٭����������3ɺ   �������Q�2������l�����l�����h����M�������\����E��u�ٝP����M�-������W�����D�����\��� ��  ���]�j h8N�������
����E�������P��\����I�����!�����x����E� �������I�����x��� ��   ǅ8���    ���8�������8���ۅ8����E��X.������AuS�E�؅P����]�M�v���������Pj Q�E��$�������P���P�M�Q���P��\����������8����M����j h(N�������3����E�������P��\����r�����J����������E� �������r��������� ��   ǅ,���    ���,�������,���ۅ,����E��X.������AuV�E�؅P����]�M�����������Pj Q�E��$�������y���P�M�z���P��\���� �����,�����t������j hN�������Y����E�������P��\���������p����������E� ���������������� ��   ǅ ���    ��� ������� ���ۅ ����E��X.������AuV�E�؅P����]�M������������Pj Q�E��$���������P�M����P��\����&����� �����h�����냋�\���������\����M���ǅ���   ǅ���    �������������ۅ����E��X.������A��  j h\N�� ����(����E�	j h ��P��������E�
j h ������������E���������� ���Pj0j j�j��������h���Q���$��8���P�y������������������������E�������R��P���Pj0j j�j��������t���Q���$��h���P�+������������������������E�������R������Pj0j j�j�������U�Q���$������P���������|�����|�����x����E���x���R������P��������t�����t�����p����E���p���R������P���������l�����l�����h����E���h���R������P��������d�����d�����`����E���`���R������P��������\�����\�����X����E���X���RV�[�������T����M������E������������E������������E������������E��������t����E��������e����E���h����V����E���8����G����E�
�������8����E�	��P����)����E� �� ��������������������u.����� t%���̉����j h �x����������M� ���� ����M��������̉����j hN�F����������M������E���(�����(���Q�<�������t�����4�����4���Q�!�������h�����@�����@���Q������j h�M��X���������E�j h�M��p���������E�����L�����X���P�MQ��p���R������P�������������������������E�������RV�z������������M�����E�������������E���p��������E� ��X�������j h�M�����������E�j h�M�������	����E�j h�M������������E����􉥠���������P�MQ������R�EP������Q������R��������������������������E�������Q�����R�������������������������E�������Q��$���R�n�������|�����|�����x����E���x���QV�H�������t����M������E���$��������E�����������E��������p����E��������a����E��������R����E� �������C����E������M�4���R��P����'���XZ�M�d�    Y_^[�Ĭ  ;�������]Ð   ������   ٻ����   ջ����   ϻ����   Ļ_$ArrayPad dauer max min �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��N����Au	��N�]�E��N����z	��N�]�E��N��N���$�f������E���E���N�X�E�_^[���   ;��Z�����]� ����������������������������������������������������U����   SVW��@����0   ��������E�$�������_^[���   ;��������]������������������������������U����   SVWQ��0����4   ������Y�M��E��@��.����Dz����E�� �M��qٝ0���م0���_^[��]�������������������������U����   SVW��8����2   ������E�@�M�Iٝ<���م<���Q�$�U��E�H�M��U�J��ٝ8���م8���Q�$�M������E_^[���   ;��������]������������������������������������������������U����   SVWQ�� ����8   ������Y�M��E��.����uǅ$���   �
ǅ$���    �E��.����uǅ ���   �
ǅ ���    ��$���3�;� ������M��E��.����z�E��ٝ$����	�Eٝ$���م$�����N���$��������E���E��.����z�E��ٝ$����	�Eٝ$���م$�����N���$�������E��X�}� u�E�� ���M���M������E�_^[���   ;��e�����]� �����������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��j��������_^[���   ;�������]� ��������������������U����   SVWQ��4����3   ������Y�M���j �EP�M�Q��c�B�H �у�;��Y���_^[���   ;��I�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���c���   ��M��B(��;������_^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��c���   �M����   ��;��b���_^[���   ;��R�����]� ����������������������������U��j�h�d�    P��  SVW��H����k  ������XD3�P�E�d�    �E�    ���]����]��E�   �M������������]ȍE�P�M�����E�P�M�
����E�P�M�Q�U�R�������M�聽���]��E��u��]�j hXO�������u����E�j h  �������_����E����􉥠���������P�MQ������R������P�=������������������������E�������RV�������������M�����E��������]����E��������N����E� �������?������̉�����j hLO�����������M�_����M�_���ǅt���    ���t�������t���ۅt����E��X.������A��   ۅt����E��u����u��]�j h\N������D����E����� ��������Pj0j j�j�Q�E��$��$���Q��������������������������E�������PV��������������M�����E���$����>����E� ������/�����t�����   ����u%���̉�<���j h �����������M�=���������M��������̉�H���j hDO�c����������M�������̉�T���j hHN�>����������M������M�����ǅh���    ���h�������h���ۅh����E��X.������A��  �E��E��]�j Q�E��$��`�������P�M�7���jj j �M������H���P�M������H�����\�����\���� �5H.ٝ����م����Q�$�h�����ٝ<�����\���� �5H.ٝ����م����Q�$������ٝ�����\����@���5H.ٝ����م����Q�$������ٝ0�����\����@���5H.ٝ����م����Q�$�R�����ٝ�����\����@�5H.ٝ����م����Q�$������ٝ$�����\����@�5H.ٝ����م����Q�$�������ٝ ���م<���؍0���ٝ����م���؍���ٝ����م����؍$���م����؍ �����ٝ����م����؍ ���م����؍$�����ٝ����م���؍0���؍$���م<���؍���؍ �����ٝ����م<���؍���؍$���م���؍0���؍ �����ٝ����Qم�����$�|������H.ٝ����م����؍����م����؍������م����؍������ٝ����م�����8O����z��ٝ������ٝ����م����ٝ�����NQم�����$������ٝ����م����ص����ٝ����م����ص����ٝ����م����ص����ٝ����j h�+��|���������E�j h ������������E�j h ������������E�j h ����������E�	����p�����|���Pj0j j�j�Qم�����$������Q�=������������������������E�
������P������Qj0j j�j�م������Q�$������R��������������������������E�������Q������Rj0j j�j�م������Q�$������P�������������������������E�������R�����Pj0j j�j�Qم�����$��$���Q�j�������������������|����E���|���P��<���Q��������x�����x�����t����E���t���P��T���Q�c�������p�����p�����l����E���l���P��l���Q�7�������h�����h�����d����E���d���P������Q��������`�����`�����\����E���\���P������Q���������X�����X�����T����E���T���P������Q��������P�����P�����L����E���L���PV��������H����M�'����E�������������E�������������E������������E���l��������E���T��������E���<��������E���$����y����E��������j����E�
�������[����E�	�������L����E�������=����E��������.����E������������E� ��|���������h�����}ԅ�u.��h��� t%���̉�����j h �q����������M�����B����M�������̉�����j h,O�?����������M�����j hO�����������E�j h�M������	����E���������������P�MQ�����R�� ���P��������������������������E�������RV��������������M�[����E��� ��������E������������E� �����������j h�N��D����f����E�j h�N��\����P����E�j h�M��t����:����E�����8�����D���P�MQ��\���R�EP��t���Q������R�������������������������E�������Q������R��������������������������E�������Q������R�������������������������E�������QV�������������M�)����E�������������E�������������E������������E���t��������E���\��������E� ��D��������E������M�{���R��P�D��n���XZ�M�d�    Y_^[�ĸ  ;��������]�   L�����   ������   ������   ��H���   ������   ��_$ArrayPad $S1 dauer max min �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������Q�E�$�������_^[���   ;�������]��������������������������������U����   SVW��<����1   �������E���$�%�����ٝ<���م<���_^[���   ;�������]����������������������������������U����   SVW��@����0   ������Q�E�$�������_^[���   ;��3�����]��������������������������������U����   SVW��<����1   �������E���$�������ٝ<���م<���_^[���   ;��������]����������������������������������U����   SVW��@����0   ������Q�E�$�}�����_^[���   ;��c�����]��������������������������������U����   SVW��<����1   �������E���$������ٝ<���م<���_^[���   ;��������]����������������������������������U����   SVW��@����0   ������Q�E�$������_^[���   ;�蓿����]��������������������������������U����   SVW��<����1   �������E���$�` ��ٝ<���م<���_^[���   ;��%�����]����������������������������������U����   SVWQ�� ����8   ������Y�M���E�P��$���Q��c�BH�H8�у�;�踾���U��
�H�J�@�B�E_^[���   ;�蒾����]� ��������������������������������������������U��j�h��d�    P���  SVW��0����q   ������XD3�P�E�d�    �E�P�M�������6����E�P�M��������V����E�P�M�Q�U�R��������M��ͩ���]����̉�H���j h �ź����@����M�m������̉�T���j h�O蠺����@����M�H������̉�`���j h�O�{�����@����M�#������̉�l���j h�O�V�����@����M�����j h �������6����E�    j h�O�����������E�����x���������Pj0j j�j�Q�E��$������Q��������@�����@�����<����E���<���P������Q������R���������8�����8�����4����E���4���QV��������0����M�8����E�������������E�������������E� ������������E������������������̉�����j h�O�,�����@����M�Է�����̉�����j h�O������@����M请���   R��P�\��X���XZ�M�d�    Y_^[���  ;��ʻ����]Ë�   d�����   ������   ������   ��dauer max min ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��0����4   ��������̉�8���j hP虷����0����M�A���_^[���   ;��}�����]��������������������������U����   SVW��$����7   ������E<P���̉�,���Q�M<������$����UR�������E<P�MQ�<������M�������=�����t�E<P�MQ�j������E<P�MQ�,������M<������脵���E��}� t<�M�����='  u �E<P�MQ�Q������E<P�MQ�H������M������E�뾋M������趢����t�E<P�MQ�������EP�������_^[���   ;��B�����]�������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���c���   ��M��B(��;�豸��_^[���   ;�衸����]������������������������������U��j�h��d�    P��$  SVW��������   ������XD3�P�E�d�    �M�����j h�P������'����E�    j h�P��L��������E�������������P��4���Q�M���������������������E������P��L���Q��d���R��������� ����� ����������E�������QV�������������M�8����E���d���������E���4���������E� ��L���������E���������������M��������̉�|���j h�P�$���������M�̲���E�   j hhP������������E�   j hXP�����������E����􉥈���������P������Q�M��������������������E������P������Q������R�������� ����� ����������E�������QV�t������������M�����E������������E������������E������������E����������������M��������̉�����j hLP�����������M袱���M�[����E�    �	�E����E��M胟��9E���  �}� u�M�*���j h�+�����衲���E�   j h ��<���舲���E�	j h ��l����r����E�
���� ��������Pj0j j�j��M�&����M�k�Q��$��$���R�����������������������E������Q��<���Rj0j j�j��M�ֹ���M�k�Q�D�$��T���R�������� ����� ����������E�������Q��l���Rj0j j�j��M腹���M�k�Q�D�$������R�K������������������������E�������Q������R�p������������������������E�������Q������R�D������������������������E�������Q������R�������������������������E�������Q������R��������������������������E�������QV��������������M�`����E������������E�������������E�������������E�������������E�������������E���T���������E�
��$��������E�	��l��������E���<��������E���������������M�����E���}��u+�}� t%���̉�����j h ����������M艮��������M�=������̉����j hXN误��������M�W����M�������̉����j h� 肯��������M�*����M�d�    Y_^[��0  ;��[�����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h�d�    P��  SVW��d�����   ������XD3�P�E�d�    ���̉�����j h�P�j����������M�����E�    �	�E���E�M����9E��(  �M�d������}����M�T����M����T>;T��  j h�P������������E�    j h�+����������E�j h�+��4����̬���E���������������P�M�����M����TR������P�x������������������������E�������R�����P�M蛺���M����TR�����P�2������������������������E�������R��4���P�M�U����M����R��L���P��������������������������E�������R��d���P��������������������������E�������R��|���P�������������������������E�������R������P�������������������������E�������R������P�g������������������������E�	������RV�A�������|����M�۩���E������������E��������x����E���|����i����E���d����Z����E���L����K����E�������<����E��������-����E���4��������E� ����������E�����������������q  j h�P�������u����E�
   j h�+�� ����\����E�j h�+��0����F����E�j h�+��`����0����E���������������P�M�E����M����TR������P��������������������������E�������R�� ���P�M������M����TR�����P�������������������������E�������R��0���P�M蹷���M����TR��H���P�P������������������������E�������R��`���P�M�s����M����R��x���P�������������������������E�������R������P�	������������������������E�������R������P��������������������������E�������R������P�������������������������E�������R������P��������|�����|�����x����E���x���R������P�Y�������t�����t�����p����E���p���R�����P�-�������l�����l�����h����E���h���RV��������d����M衦���E�������M����E��������>����E��������/����E�������� ����E������������E������������E���x���������E���H���������E������������E�������������E���`��������E���0��������E�
�� ��������E����������������������̉� ���j h� ������������M袥���M�d�    Y_^[�Ĝ  ;��ө����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h\�d�    P��  SVW��L�����   ������XD3�P�E�d�    �E�    �M�������{����E��}� t#�M������=�  u�E�   �M��)����E��׃}� uj h�  �M蝩����蔡���E�   �M臩���������E��}� �s  �M�蛰��=�  �P  �M�X������]����E��E�    ���̉�����j hQ�����������M赢�����̉�����j h�P�����������M萢���M萳�����̉�����j h�P軣���������M�c����M�c����E�    �	�E����E��M�����9E��/  �M譱�����}����M蝱���M����T>;T�  �E�    �	�E����E��}���  �}� u�M����j h�+�����������E�    j h �����������E�j h ����������E����􉥰���������Pj0j j�j��M�k��U�Q�
�$������P�k������������������������E�������R������Pj0j j�j��M�k��U�Q�D
�$�����P��������|�����|�����x����E���x���R�����Pj0j j�j��M�k��U�Q�D
�$��4���P�Ӻ������t�����t�����p����E���p���R��L���P���������l�����l�����h����E���h���R��d���P�̹������d�����d�����`����E���`���R��|���P蠹������\�����\�����X����E���X���R������P�t�������T�����T�����P����E�	��P���RV�N�������L����M�����E�������蔼���E���|���腼���E���d����v����E���L����g����E���4����X����E�������I����E��������:����E�������+����E� �����������E������������
����M�����E����E��6����E����E����̉�����j h �c����������M������  �E�    �	�E����E��}���  �}� u�M蝿��j h�+�����������E�
   j h ������������E�j h ��$��������E����􉥸���������Pj0j j�j��M�k��U�Q�
�$������P�e������������������������E�������R������Pj0j j�j��M�k��U�Q�D
�$�����P��������|�����|�����x����E���x���R��$���Pj0j j�j��M�k��U�Q�D
�$��<���P�ͷ������t�����t�����p����E���p���R��T���P��������l�����l�����h����E���h���R��l���P�ƶ������d�����d�����`����E���`���R������P蚶������\�����\�����X����E���X���R������P�n�������T�����T�����P����E���P���RV�H�������L����M�����E�������莹���E������������E���l����p����E���T����a����E���<����R����E�������C����E��������4����E���$����%����E�
�����������E����������������M�����E����E��6������̉�����j h �f����������M�����������̉�����j h� �<����������M�����M�����M�������̉�����j h� �����������M诛���E�P�a������M��z����E������}� uj h�  �M����������R��P����%���XZ�M�d�    Y_^[�Ĵ  ;�藟����]ÍI    ������   ��phongNormal ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P��  SVW��������  ������XD3�P�E�d�    �M������E�    �E�    �E�    �M�������蕘���E��}� �u  �M�����='  �:  �E����E��E؃��E؋E��E�j htQ������苙���E�    j hhQ�������r����E�j hXQ�� ����\����E����􉥔���������P�M�Q������R�������������������������E�������Q������R������P�M������������������������E�������R�� ���P�����Q�۰������|�����|�����x����E���x���P��0���Q诰������t�����t�����p����E���p���P��H���Q胰������l�����l�����h����E���h���PV�]�������d����M������E���H���裳���E���0���蔳���E������腳���E��������v����E��������g����E��� ����X����E� �������I����E������������7����M�|������̉�`���j hLQ觗���������M�O����E�    �	�E����E��M����9E���  �E�P��d���Q�M��j����M莥�����}����M�~����M����T>;T�F  Qمl����$Qمh����$Qمd����$��P����6���Qمx����$Qمt����$Qمp����$��<�������Q�E��$Q�E��$Qم|����$��(�������Q�E��$Q�E��$Q�E��$������ʾ��Q�HQ�$Q���$Q���$��l���詾��PQ���$Q�HQ�$Q���$������臾��PQ���$Q���$Q���$�������i���P������P�M�T����������P�������]�����P���P������Q������R衲�������P����P��T����@��X�����<���P������Q������R�j��������<����P��@����@��D�����(���P������Q������R�3��������(����P��,����@��0��������P������Q������R��������������P������@�����j hDQ������0����E�   j h ��H��������E�	j h�+��x��������E�
j h �����������E�j h�+�������Ք���E�j h �����返���E�������������Pj0j j�j�Qم,����$��0���Q�E������������������������E�������P��H���Qj0j j�j�Qم(����$��`���R� ������������������������E�������Q��x���Rj0j j�j�Qم@����$������P軬������|�����|�����x����E���x���R������Pj0j j�j�Qم<����$������Q�v�������t�����t�����p����E���p���P������Qj0j j�j�QمT����$������R�1�������l�����l�����h����E���h���Q�����Rj0j j�j�QمP����$�� ���P��������d�����d�����`����E���`���R��8���P��������\�����\�����X����E���X���R��P���P��������T�����T�����P����E���P���R��h���P蹪������L�����L�����H����E���H���R������P荪������D�����D�����@����E���@���R������P�a�������<�����<�����8����E���8���R������P�5�������4�����4�����0����E���0���R������P�	�������,�����,�����(����E���(���R������P�ݩ������$�����$����� ����E��� ���R������P豩��������������������E������R�����P腩��������������������E������RV�_�����������M������E������襬���E�������薬���E�������臬���E��������x����E��������i����E��������Z����E��������K����E���h����<����E���P����-����E���8��������E��� ��������E�������� ����E������������E������������E���`����ӫ���E���0����ī���E������赫���E�������覫���E�
������藫���E�	��x���舫���E���H����y����E�����������g����	  Qمl����$Qمh����$Qمd����$����������Qمx����$Qمt����$Qمp����$�������Ƿ��Q�E��$Q�E��$Qم|����$������褷��Q�E��$Q�E��$Q�E��$������脷��Q�HQ�$Q���$Q���$��(����c���PQ���$Q�HQ�$Q���$��<����A���PQ���$Q���$Q���$��P����#���P��d���P�M������贠��P��T�������������P��T���Q��x���R�[�������������P�������@������������P��T���Q������R�$�������������P�������@������������P��T���Q������R��������������P�������@������������P��T���Q������R趪������������P�������@������j hDQ�����������E�   j h ������э���E�j h�+��4���軍���E� j h ��d���襍���E�!j h�+������菍���E�"j h �������y����E�#j h�+�������c����E�$j h ��$����M����E�%��������������Pj0j j�j�Qم�����$������Q�ӥ�����������������������E�&������P�����Qj0j j�j�Qم�����$�����R莥�����������������������E�'������Q��4���Rj0j j�j�Qم�����$��L���P�I�������|�����|�����x����E�(��x���R��d���Pj0j j�j�Qم�����$��|���Q��������t�����t�����p����E�)��p���P������Qj0j j�j�Qم�����$������R迤������l�����l�����h����E�*��h���Q������Rj0j j�j�Qم�����$������P�z�������d�����d�����`����E�+��`���R������Pj0j j�j�Qم�����$�����Q�5�������\�����\�����X����E�,��X���P��$���Qj0j j�j�Qم�����$��<���R��������T�����T�����P����E�-��P���Q��T���R��������L�����L�����H����E�.��H���Q��l���R��������D�����D�����@����E�/��@���Q������R轢������<�����<�����8����E�0��8���Q������R葢������4�����4�����0����E�1��0���Q������R�e�������,�����,�����(����E�2��(���Q������R�9�������$�����$����� ����E�3�� ���Q������R����������������������E�4�����Q������R����������������������E�5�����Q�����R赡��������������������E�6�����Q��,���R艡���������������� ����E�7�� ���Q��D���R�]������������������������E�8������Q��\���R�1������������������������E�9������Q��t���R�������������������������E�:������Q������R�٠�����������������������E�;������QV賠�����������M�M����E�:������������E�9��t��������E�8��\����ۣ���E�7��D����̣���E�6��,���轣���E�5�����讣���E�4������蟣���E�3������萣���E�2������聣���E�1�������r����E�0�������c����E�/�������T����E�.��l����E����E�-��T����6����E�,��<����'����E�+����������E�*�������	����E�)������������E�(��|��������E�'��L����ܢ���E�&������͢���E�%������辢���E�$��$���询���E�#������蠢���E�"������葢���E�!������肢���E� ��d����s����E���4����d����E�������U����E������������C����=������̉�����j hXN趆���������M�^����M�	������̉�����j h� 艆���������M�1����M��ƒ��=�  u	�E����E��M�������E������E�    �}��	  ǅH���   ���H�������H�����H���;E���  j h4Q�����������E�<   j h,Q�����������E�=j h Q��(����ׅ���E�>���􉥼���������P������Q�M詘���������������������E�?������P������Q��H���R�����P�\������������������������E�@������R��(���P��@���Q�S�������|�����|�����x����E�A��x���P��X���Q�'�������t�����t�����p����E�B��p���P��p���Q���������l�����l�����h����E�C��h���PV�՜������d����M�o����E�B��p��������E�A��X��������E�@��@���������E�?����������E�>�������ߟ���E�=��(����П���E�<������������E�����������诟������R��P�	�z��XZ�M�d�    Y_^[��$  ;�������]ÍI     	����   �	d���0   �	P���   �	<���   �	(���   �	���   �	����0   �	����   �	����   �	����   �	����   �	T���0   �	mirrorX d c b a mirrorX d c b a uvwKoord texturCoord �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��/����M����$����M��������M���$�����E�M����P�Q�@�A�E�M������P�Q�@�A�E�M������P�Q�@�A�E�M���$���P�Q�@�A�E�_^[���   ;������]� ����������������������������������������������������������U����   SVW��4����3   ������E�@�M�	�U�B�E�@ �M�I���U�B,�E�H��ٝ<���م<���Q�$�M�A�U�
�E�@�M�A�U�J���E�@(�M�I��ٝ8���م8���Q�$�U�B�E��M��U�B�E�H���M�A$�U�J��ٝ4���م4���Q�$�M躣���E_^[���   ;��~����]��������������������������������������������������������������U���  SVWQ�������A   ������Y�M��M��n����E�P�MQ�U�R��c�HD�Q<�҃�;���}���   �u��}�ER��P�h	�Bq��XZ_^[��  ;��}����]� �   p	����0   |	us �������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��/����M����$����M��������M���$�����E�_^[���   ;��}����]������������������������������U��j�h��d�    P��  SVW��`����%  ������XD3�P�E�d�    �E�    �M��~�����[x���E��}� t%�M��݅��=�  u	�E���E�M��v���E����E�    �}� u*���̉�����j h�Q�Iy���������M��w����   j h�Q�������$y���E�    j h�Q������y���E���������������P�Mԃ�Q������R�Ü�����������������������E�������Q�����R�� ���P躐�����������������������E�������RV蔐�����������M�.w���E��� ����ړ���E��������˓���E� �����輓���E�����������誓���E�    �E�    �	�E����E��M����9E���  �M�:������}����M�*����M����T>;T��  j h�Q��D�����w���E�   j h�+��t����w���E�j h�+�������w���E�j h �������w���E�����8�����D���P�Mȃ�Q��\���R�D������������������������E�������Q��t���R�Eȃ�P������Q�
������������������������E�	������P������Q�U�R������P�Ӛ�����������������������E�
������R������P������Q�ʎ�����������������������E�������P�����Q螎�����������������������E�������P�����Q�r������������������������E�������P��4���Q�F������������������������E�������P��L���Q��������������������|����E���|���PV��������x����M�t���E���L����:����E���4����+����E�����������E�����������E�
������������E�	�����������E�������������E���\����ѐ���E�����������E�������賐���E���t���褐���E�������D���蒐���Eȃ��E��  j h�Q��p����u���E�   j h�+��������t���E�j h�+��������t���E�j h�+�� ����t���E�j h ��0����t���E�����d�����p���P�Mȃ�Q������R�^������������������������E�������Q������R�Eȃ�P������Q�$������������������������E�������P������Q�Uȃ�R������P�������������������������E�������R�� ���P�M�Q�����R賗�����������������������E�������Q��0���R��H���P誋�����������������������E�������R��`���P�~������������������������E�������R��x���P�R������������������������E�������R������P�&�������������������|����E���|���R������P���������x�����x�����t����E���t���R������P�Ί������p�����p�����l����E���l���R������P袊������h�����h�����d����E���d���RV�|�������`����M�q���E�����������E�������賍���E�������褍���E�������蕍���E���x���膍���E���`����w����E���H����h����E�������Y����E��������J����E��������;����E��������,����E���0��������E��� ��������E�������������E�������������E�������p����ތ���Eȃ��E��6������̉�����j hXN�Hq���������M��o���Eԃ��EԋE�;E�������M�d�    Y_^[�Ġ  ;��t����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hx�d�    P��  SVW��@�����   ������XD3�P�E�d�    �E�    �M�s�����+m���E��}� t#�M��z��=�  u�E�   �M���j���E��׃}� uj h�  �M�Ms�����Dk���M�>s������l���E��}� �y  �M��Rz��=�  �V  ���̉�����j h�Q��m���������M�l���E�    �E�    �	�Eȃ��EȋM����9E���  �M��{�����}����M��{���M����T>;T�i  j h�P�������gm���E�    j h�+�������Nm���E�j h�+������8m���E����􉥤���������P�Mԃ�Q������R�������������������������E�������Q������R�Eԃ�P������Q趐�����������������������E�������P�����Q�U�R��(���P��������������������|����E���|���R��@���P�}�������x�����x�����t����E���t���R��X���P�Q�������p�����p�����l����E���l���R��p���P�%�������h�����h�����d����E���d���R������P���������`�����`�����\����E�	��\���RV�Ӄ������X����M�mj���E������������E���p����
����E���X���������E���@��������E���(����݆���E��������Ά���E�������迆���E������谆���E� ������衆���E�����������菆���Eԃ��E��H  j h�P��������j���E�
   j h�+��������j���E�j h�+�������j���E�j h�+��<����j���E����􉥠���������P�Mԃ�Q������R�q������������������������E�������Q������R�Eԃ�P������Q�7������������������������E�������P�����Q�Uԃ�R��$���P���������������������|����E���|���R��<���P�M�Q��T���R�ƍ������x�����x�����t����E���t���Q��l���R�ā������p�����p�����l����E���l���Q������R蘁������h�����h�����d����E���d���Q������R�l�������`�����`�����\����E���\���Q������R�@�������X�����X�����T����E���T���Q������R��������P�����P�����L����E���L���Q������R��������H�����H�����D����E���D���QV�������@����M�\g���E������������E�������������E������������E��������ۃ���E��������̃���E���l���轃���E���T���讃���E���$���蟃���E�������萃���E�������聃���E���<����r����E�������c����E�
�������T����E������������B����Eԃ��E��������̉�����j h� �g���������M�Tf���M��+d���E��}����}� uj h�  �M�l�����n���M�d�    Y_^[���  ;��Yj����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P���
  SVW��4�����  ������XD3ŉE�P�E�d�    �E�    j h�S�������e���E�j h  ��������d���E�����|���������P�MQ������R������P��|������t�����t�����p����E���p���RV�|������l����M�Qc���E������������E������������E� �����������M�$t���E�    �E�    �M��<n�����]�j hL�M��<d���E��M��n�����]���ٝx�����ٝl�����ٝ`�����H����Ho���E�ǅ<���    �M�i�����b����0�����0��� �(  ��0���� p��=�  ��  ��0�����$���j ��$����x�������������<������������� ��  j hL�������sc���E�������P��H���螁���E��������~��ǅ ���    ��� ������� ����� ����C  ǅ����    ������do��=G  u�����������Q���$Q���$Q���$�������	�����M��P�U��@�E����]������� ��  �� ���P�������aq������  �� �����t�����t��� t��t����/  ��t����q  �  �������Ql��Ph4  �����P������Ӌ����MȋP�Ű@�E�Q���$h5  ������Ja���]��� ���P�����蝀���E܍�@����Cm����t�����t�����p����E���p���Qh�  ��X���R��$���P�M���f����l�����l�����h����E���h����n����d�����d�����`����E�	��`���P��H��������E���X�����|���E���$����T���E���@�����|���k��p����4k��Ph`	  ������P�����越����M��P�U��@�E�Q���$ha	  ������-`���]��Q���$h�  ������`��ٝx��������Eȉ������M̉������UЉ�����j hL�������`���E�
������P��H����Fe���������E���������{�������� tJ�M萋����������t7Q���$Q���$Q���$�������z�����������P�������@������مx�����S�xS�5hSٝl���مl���ٝ�����E�ٝ�����E�ٝ�����E�ٝ����م�����XSم�����HS��م�����8S��ٝ����م�����M�����ٝ`����M���������p��ٝ������<��� ��
  ������ڂ�������������̉�����P�mo����t���V�]������p�����p�����l����M����j h$S�������._���E�j hS��0����_���E���������������P������L������̉����P��n����t��������Q��\������p�����p�����l����E���l���P��0���Q��H���R�v������h�����h�����d����E���d���QV�v������`����M� ]���E���H�����y���E�������y���E���0����y���E��������y���M��m�����̉�`���j h�R�^����t����M�\���M�m��j h�R��x�����]���E�j h�R��������]���E�����l�����x���Pj0j j�j�Qم�����$������Q�Wv������t�����t�����p����E���p���P������Q������R�uu������l�����l�����h����E���h���QV�Ou������d����M��[���E��������x���E��������x���E��������wx���E���x����hx��j h ��������\���E�j h �������\���E�j h ��D����\���E�j h�R��t����\���E���������������Pj0j j�j�Qم�����$������Q�)u������t�����t�����p����E���p���P�����Qj0j j�j�Qم�����$��,���R��t������l�����l�����h����E���h���Q��D���Rj0j j�j�Qم�����$��\���P�t������d�����d�����`����E���`���R��t���P������Q�s������\�����\�����X����E���X���P������Q�s������T�����T�����P����E���P���P������Q�es������L�����L�����H����E���H���P������Q�9s������D�����D�����@����E���@���P������Q�s������<�����<�����8����E���8���PV��r������4����M�Y���E��������-v���E��������v���E��������v���E�������� v���E���������u���E���\�����u���E���,�����u���E���������u���E���t����u���E���D����u���E�������u���E��������u��j h ������Z���E�j h ��@�����Y���E� j h ��p�����Y���E�!j h�R��������Y���E�"������������Pj0j j�j�Qم�����$��(���Q�Ir������t�����t�����p����E�#��p���P��@���Qj0j j�j�Qم�����$��X���R�r������l�����l�����h����E�$��h���Q��p���Rj0j j�j�Qم�����$������P�q������d�����d�����`����E�%��`���R������P������Q��p������\�����\�����X����E�&��X���P������Q�p������T�����T�����P����E�'��P���P������Q�p������L�����L�����H����E�(��H���P�� ���Q�Yp������D�����D�����@����E�)��@���P�����Q�-p������<�����<�����8����E�*��8���PV�p������4����M�V���E�)������Ms���E�(�� ����>s���E�'�������/s���E�&������� s���E�%�������s���E�$�������s���E�#��X�����r���E�"��(�����r���E�!��������r���E� ��p�����r���E���@����r���E�������r��j h ��<����%W���E�+j h�R��l����W���E�,����0�����<���Pj0j j�j�Qمl����$��T���Q�o������t�����t�����p����E�-��p���P��l���Q������R�n������l�����l�����h����E�.��h���QV�n������d����M�'U���E�-��������q���E�,��T�����q���E�+��l����q���E���<����q��j h �������#V���E�/j h�R�������V���E�0���􉥜���������Pj0j j�j�Qم`����$������Q�n������t�����t�����p����E�1��p���P������Q������R�m������l�����l�����h����E�2��h���QV�m������d����M�%T���E�1��������p���E�0��������p���E�/�������p���E��������p���M�x�����̉����j h�R�U����t����M�S��j hL�� �����T���E�3�� ���P��H����Y��������E��� ����:p������� ��  ������P�M�`j����t�����t�����p����E�4��p���R���̉�D�����H���P�}d����l�����P���Q�	q������h�����h�����d����E�5��d���P��x���Q�M�5W����`�����`�����\����E�6��\����Y����;����E�5��x����W���E�4��P�����U���E��������W����;������  j h ��������S���E�7j htR�������S���E�8���􉥠���������P���̉�������H���R�c����t���������P�Q������p�����p�����l����E�9��l���R������P�� ���Q�Fk������h�����h�����d����E�:��d���PV� k������`����M�Q���E�9�� ����fn���E�8�������Wn���E�7�������Hn���E��������9n����  j hTR��$����R���E�;j h8R��`����R���E�<���������H���P��$���Q���̉�<�����H���R�kb����t�����H���P�P������p�����p�����l����E�=��l���R��`���P��x���Q�-j������h�����h�����d����E�>��d���P������Q�j������`�����`�����\����E�?��\���PV��i������X����M�uP���E�>�������!m���E�=��x����m���E�<��H����m���E�;��`�����l���E���$�����l���M��p�����̉�����j h0R�UQ����t����M��O�����̉�������H���P�4a����t���������Q��m������p�����p�����l����E�@��l���P������Q�M�(E����������G���E���������R����<�������<�����0����PM����0����������<��� t-�M�t�����̉� ���j h� �P����t����M�0O����<��� ��  j hL��0����[P���E�A��0���P�����Q�M��<����t�����t�����p����E�B��p�����T��������E�A������|k���E���0����mk������� ��   j h ��T�����O���E�Cj hR��������O���E�D����H�����T���P��l���Q�M�3<����t�����t�����p����E�E��p���P������Q������R�}g������l�����l�����h����E�F��h���QV�Wg������d����M��M���E�E�������j���E�D��l����j���E�C�������j���E���T����pj���   ���̉�����j h�Q��N����t����M�M���M�^�����̉�����j h�Q�N����t����M�^M���M�	r���M�r�����̉�����j h� �N����t����M�)M���E���H�����i���E� �M���i���E������M�i��R��P�F	�D��XZ�M�d�    Y_^[�M�3��f�����
  ;��Q����]Ð   F	����   �F	����   ~F	����   lF	H���   aF	����   TF	diffuseColor texturName TransparencyColor ColorTexName ColorColor ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M���8�������_^[���   ;��KJ����]� ���������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BT�H,�у�;���I��_^[���   ;���I����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BT�H0�у�;��kI��_^[���   ;��[I����]� �������������������������������������U����   SVW��$����7   ������M�qi�����̉�,���j h� ��E����$����M�D���M�Di���M�<i�����̉�8���j h� �E����$����M�dD��_^[���   ;��H����]����������������������������������������%T�U����   SVW��<����1   ������} t�E��<������c�x4����<�����<���Q�UR�EP��l����_^[���   ;��
H����]���������������������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��M��Sg��_^[���   ;���F����]������������������U����   SVWQ������:   ������Y�M��E��x t�   �E��8 t)��E��Q��c�B<�H�у�;��F���E��     �E��x tS�E��x t@�E��H��,�����,����� ����� ��� tj�� ����jj��������
ǅ���    �E��@    _^[���   ;��F����]���������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��B:���E��t�E�P�bY�����E�_^[���   ;��~E����]� ������������������������U����   SVWQ������?   ������Y�M������P��c����P�M��d�������������9�������_^[���   ;���D����]���������������������������U����   SVWQ��$����7   ������Y�M��E��x ufh�S�@B��Phij�5������,�����,��� t�MQ��,����R����$����
ǅ$���    �U���$����B�E��x u3��Q�E��x t�E�3Ƀ8 �����9��EP��c�Q<��Ѓ�;��D���M���E��@   �E�3Ƀ8 ����_^[���   ;���C����]� �����������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@   ��c�H<��Q��;��]C���M���E�3Ƀ8 ����_^[���   ;��;C����]����������������������������������������U����   SVWQ��4����3   ������Y�M��E��x t�   �O�E��x u3��B��E��Q��c�B<�H�у�;��B���E��     �E��@    �E��HQ�M��ja��_^[���   ;��~B����]�������������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 u��c�H��#��EP�M��R��c�H<�Q�҃�;���A��_^[���   ;���A����]� ��������������������������������U����   SVW��@����0   �����󫹔c��a��_^[���   ;��A����]���������������������U����   SVW��@����0   ������EP��c�yW��_^[���   ;��4A����]�����������������U���  SVW�������C   ������XD3ŉE��EP��c�W��P�M���M��j h�S�������=��j �E�P�����Q�M��lH�������������������Y����������t�M��H���M���X���E�5j�E�P�M���8���EP�M�Q�M���[���E�P�M�ZM���M��X���ER��P�W	�3��XZ_^[�M�3��U����  ;��"@����]Ë�   W	����   (W	����   $W	str pos ������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q�B$�Ѓ�;��S?��_^[���   ;��C?����]� �����������������������������U���0  SVW�������L   ������XD3ŉE��EP��c�U��P�M���K��j h�S��������;��j �E�P������Q�M��lF��������������������W����������t�M��F���M���V���E�   j�E�P�M���6���EP�M�Q�M���Y��j h�S������M;��j �E�P�����Q�M���E�������������������V����������t�M�MF���M��vV���E�5j�E�P�M��j6���EP�M�Q�M��UY���E�P�M��J���M��?V���ER��P��Y	�/1��XZ_^[�M�3��S����0  ;��=����]Ë�   �Y	����   �Y	����   �Y	str pos ��������������������������������������������������������������������������������������������������������������������U���T  SVW�������U   ������XD3ŉE��EP��c��R��P�M���I��j h�S�������9��j �E�P������Q�M��LD���������������������T����������t�M�D���M���T���E�2  j�E�P�M���4���EP�M�Q�M��W��j h�S�������-9��j �E�P������Q�M���C��������������������qT����������t�M�-D���M��VT���E�   j�E�P�M��G4���EP�M�Q�M��2W��j h�S������8��j �E�P�����Q�M��LC��������������������S����������t�M�C���M���S���E�5j�E�P�M���3���EP�M�Q�M��V���E�P�M�:H���M��S���ER��P�$\	�.��XZ_^[�M�3��|P����T  ;��;����]Ë�   ,\	����   H\	����   D\	str pos ����������������������������������������������������������������������������������������������������������������������������������������������������U���x  SVW�������^   ������XD3ŉE��EP��c�?P��P�M��G��j h�S��������6��j �E�P������Q�M��A��������������������1R����������t�M��A���M��R���E�  j�E�P�M��2���EP�M�Q�M���T��j h�S�������m6��j �E�P������Q�M��A��������������������Q����������t�M�mA���M��Q���E�2  j�E�P�M��1���EP�M�Q�M��rT��j h�S��������5��j �E�P������Q�M��@��������������������1Q����������t�M��@���M��Q���E�   j�E�P�M��1���EP�M�Q�M���S��j h�S������m5��j �E�P�����Q�M��@�������������������P����������t�M�m@���M��P���E�5j�E�P�M��0���EP�M�Q�M��uS���E�P�M��D���M��_P���ER��P�d_	�O+��XZ_^[�M�3��<M����x  ;���7����]Ë�   l_	����   �_	����   �_	str pos ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �������EP��c�Q<�B�Ѓ�;��6��_^[���   ;��6����]���������������������������������U���p  SVW�������\   ������ǅ����    j h T�������43��P�'�����E��������N���}� u3���   �E�    �E�P�M���+���E�P�M�Q�M��l6������   �}���   �M��D+���E��}� tF�EP��������=��������Pj������Q�M��?������������&����tǅ����   �
ǅ����    ��������������������t���������������M����������t��������������M����������t�EԉE�������E�R��P�,b	�}(��XZ_^[��p  ;���4����]Ë�   4b	����   cb	����   _b	����   Xb	browse dat id ��������������������������������������������������������������������������������������������������������������������������U����   SVW������:   ������} u3��   �EP�M���)���E�    �E�    �E�P�M�Q�M��h4����tT�}�t�}�u"�EP�M��>)��P�x*������t�   �*�$�}�u�EP�M��L������$����t�   ��3�R��P��c	��&��XZ_^[���   ;��p3����]�   �c	����   �c	����   �c	����   �c	dat id browse ����������������������������������������������������������������������������������U����   SVW��@����0   �����󫡨c�H<��Q��;��2��_^[���   ;��2����]�������������������������U����   SVW��@����0   �������j���c�H�Q�҃�;��G2��_^[���   ;��72����]��������������������U����   SVW��@����0   �������EP��c�Q�B�Ѓ�;���1��_^[���   ;���1����]���������������������������������U����   SVW��@����0   �������EP��c�Q�B�Ѓ�;��t1��_^[���   ;��d1����]���������������������������������U����   SVWQ��4����3   ������Y�M���j��E�P��c�Q���   �Ѓ�;���0���E�_^[���   ;���0����]������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B���   �у�;��x0���E�_^[���   ;��e0����]� �������������������������������U����   SVWQ��4����3   ������Y�M���j��E�P��c�Q���   �Ѓ�;���/����j �E�P�MQ��c�B���   �у�;���/���E�_^[���   ;���/����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q�B�Ѓ�;��O/��_^[���   ;��?/����]����������������������������U����   SVWQ��4����3   ������Y�M���j �E�P�MQ��c�B���   �у�;���.���E�_^[���   ;���.����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H���   �҃�;��U.��_^[���   ;��E.����]� �������������������������������U����   SVWQ��(����6   ������Y�M���j���c�H�Q�҃�;���-���E�}� u3��+��EP�M�Q�U�R��c�H���   �҃�;��-���E�_^[���   ;��-����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H�у�;��+-��_^[���   ;��-����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H�у�;��,�������_^[���   ;��,����]� ������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q�B�Ѓ�;��/,��_^[���   ;��,����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q�B�Ѓ�;��+��_^[���   ;��+����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H�у�;��K+��_^[���   ;��;+����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�Hh�у�;���*��_^[���   ;��*����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�Ht�у�;��K*��_^[���   ;��;*����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�Hl�у�;���)��_^[���   ;��)����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�Hp�у�;��K)��_^[���   ;��;)����]� �������������������������������������U����   SVWQ��(����6   ������Y�M���EP�M�Q��c�B�Hl�у�;���(���E�}��u3��"��E�P�M�Q��c�B�H|�у�;��(��_^[���   ;��(����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H|�у�;��(��_^[���   ;��(����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M���(�����u�E�"��EP�M�Q��c�B�HH�у�;��'��_^[���   ;��u'����]� �������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��4(�����u�E�"��EP�M�Q��c�B�HL�у�;���&��_^[���   ;���&����]� �������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��'�����u�E�U�%��EP�M�Q��c�B���   �у�;��_&��_^[���   ;��O&����]� �����������������������������������������U����   SVWQ��(����6   ������Y�M��EP�M��'�����u�E�B��EP�M�Q��c�B���   �у�;���%���E�M���,����u
�M���8����E_^[���   ;��%����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��D&�����u�E�"��EP�M�Q��c�B�HD�у�;��%��_^[���   ;���$����]� �������������������������������U����   SVWQ�� ����8   ������Y�M��EP�M��%�����u�E�M���P�Q�@�A�E�>��EP�M�Q��$���R��c�H�Q`�҃�;��Y$���M���P�Q�@�A�E_^[���   ;��3$����]� ���������������������������������������������U���  SVWQ�������A   ������Y�M��EP�M���$�����u�u�   �}�E�7��EP�M�Q�� ���R��c�H�Qd�҃�;��#���   ���}�E_^[��  ;��s#����]� ���������������������������������������������U����   SVWQ������=   ������Y�XD3ŉE��M�EP�M��$�����u�EP�M��/���E�b��EP�M�Q��c�B�HP�у�;���"���E�M��+���}� t�E�P�M���=���E�P��&�����E�P�M�/���M��;���ER��P��t	����XZ_^[�M�3���7�����   ;��d"����]� ��   �t	����   �t	����   �t	s str ����������������������������������������������������������������������U����   SVW��@����0   ������E�8 t ��E�Q��c�B�H�у�;��!���E�     _^[���   ;��!����]������������������������������U���   SVWQ�� ����@   ������Y�XD3ŉE��M�EP�M��J"�����u�EP�M�.���E�b��EP�M�Q��c�B�HT�у�;��� ���E�M��+���}� t�E�P�M��.���E�P�P@�����E�P�M�X.���M��_���ER��P��v	�!��XZ_^[�M�3��6����   ;�� ����]� ��   �v	����   �v	����   �v	f fn �����������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M���EP�M�Q��c�B�H\�у�;������E�}� t�E�P�M�VI���E��M�|���E_^[���   ;������]� ��������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H\�у�;��;��_^[���   ;��+����]� �������������������������������������U����   SVWQ��$����7   ������Y�M��EP�M��������u�E��P�E��P�E�8��EP�M�Q��(���R��c�H�QX�҃�;������P�E��P�E_^[���   ;��o����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H�Q$�҃�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H�Q(�҃�;��x��_^[���   ;��h����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q���   �Ѓ�;�����_^[���   ;�������]� ��������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$�EP�M�Q��c�B�H �у�;��t��_^[���   ;��d����]� ������������������������������U����   SVWQ��$����7   ������Y�M�j �EP�M��!
����E�P�MQ�U�R��c�H���   �҃�;������M��;)��R��P�h{	�A��XZ_^[���   ;������]�    p{	����   |{	data �����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H�Q<�҃�;��(��_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H�Q@�҃�;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H�Q,�҃�;��(��_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H�Q0�҃�;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H�Q8�҃�;��(��_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H�Q4�҃�;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B���   �у�;��(��_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H���   �҃�;����_^[���   ;������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q���   �Ѓ�;�� ��_^[���   ;������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H���   �҃�;����_^[���   ;������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B���   �у�;��(��_^[���   ;������]� ����������������������������������U����   SVWQ��(����6   ������Y�M��EP�M��'-���E�M���5��_^[���   ;������]� ��������������������������������U����   SVWQ��(����6   ������Y�M��EP�M��,���E�EP�MQ�M����_^[���   ;��.����]� ������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q���   �Ѓ�;�����_^[���   ;������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H���   �҃�;��E��_^[���   ;��5����]� �������������������������������U����   SVWQ��4����3   ������Y�M���h#  �EP�MQ�U�R��c�H���   �҃�;�����_^[���   ;������]� ��������������������������U����   SVWQ��4����3   ������Y�M���hF  �EP�MQ�U�R��c�H���   �҃�;��@��_^[���   ;��0����]� ��������������������������U����   SVWQ��(����6   ������Y�M��EP�M��G*���E�EP�M��*��_^[���   ;�������]� ����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B���   �у�;��X��_^[���   ;��H����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H���   �҃�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H���   �҃�;��U��_^[���   ;��E����]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E�_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��    �E��M�H�E�_^[��]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��M�H�E�_^[��]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��E�X�E�_^[��]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E�E��X�E�_^[��]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q��c���   �H�у�;������E�_^[���   ;�������]� ��������������������������������������������U����   SVWQ������:   ������Y�XD3ŉE��M�j �EP�M��s���E��     �E��@    ��E�P�M�Q��c���   �H$�у�;��=���M��&���E�R��P� �	���XZ_^[�M�3��#�����   ;������]� �   (�	����   4�	str ��������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q��c���   �H$�у�;��U���E�_^[���   ;��B����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q��c���   �H0�у�;�����E�_^[���   ;������]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q��c���   �H �у�;�����E�_^[���   ;������]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q��c���   �H(�у�;��u���E�_^[���   ;��b����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q��c���   �H,�у�;���
���E�_^[���   ;���
����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��j �EP�M�Q��c���   �H�у�;��3
���E�_^[���   ;�� 
����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q��c���   �H4�у�;��	���E�_^[���   ;��	����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��M�H�E�_^[��]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�MQ�U�R��c���   �Qh�҃�;�����E�_^[���   ;������]� �����������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�MQ�U�R��c���   �Q\�҃�;������E�_^[���   ;�������]� �����������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q��c���   �Hd�у�;��U���E�_^[���   ;��B����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c���   �H�у�;�����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c���   �H�у�;��H�������_^[���   ;��1����]� ���������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�UR��c���   �Q�҃�;�����_^[���   ;������]� �������������������������������U����   SVWQ��4����3   ������Y�M�j �E�P�M����E�_^[���   ;��L����]� ����������������������U����   SVWQ��4����3   ������Y�M���E�P��c���   ��Ѓ�;�����_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M���E�P��c���   ��Ѓ�;��}��_^[���   ;��m����]��������������������������U����   SVWQ��4����3   ������Y�M���E�P��c���   �B�Ѓ�;����_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c���   �B8�Ѓ�;����_^[���   ;������]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c���   �Bl�Ѓ�;��,��_^[���   ;������]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c���   �B<�Ѓ�;����_^[���   ;������]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c���   �B@�Ѓ�;��L��_^[���   ;��<����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c���   �BH�Ѓ�;�����_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c���   �BT�Ѓ�;��l��_^[���   ;��\����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c���   �BD�Ѓ�;��� ��_^[���   ;��� ����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c���   �BL�Ѓ�;�� ��_^[���   ;��| ����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c���   �BP�Ѓ�;�� ��_^[���   ;�� ����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c���   �BX�Ѓ�;�����_^[���   ;�������]�������������������������U����   SVWQ��(����6   ������Y�M���E�P��c���   �BX�Ѓ�;��<����E�}� u3���EP�MQ�M��(��_^[���   ;�������]� �����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c���   �Q�҃�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��(����6   ������Y�M���E�P��c���   �BX�Ѓ�;������E�}� u3���EP�MQ�M��|��_^[���   ;��������]� �����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c���   �Q8�҃�;��u���_^[���   ;��e�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���j�E�P��c���   �B`�Ѓ�;������_^[���   ;��������]�����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c���   �H`�у�;�����_^[���   ;��x�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E��M���j j j �E��Q��c�B���   �у�;�������U��B�E�_^[���   ;��������]� �����������������������������U����   SVWQ��4����3   ������Y�M���j j j �E��Q��c�B���   �у�;��t����U��B_^[���   ;��^�����]���������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��<��E��HQ�UR�EP�M��R��c�H���   �҃�;�������M��A�   _^[���   ;��������]� ����������������������������������������������U����   SVW��@����0   ������E��c��c� _^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��E��� P������_^[���   ;��������]���������������������������U����   SVW��@����0   �������EP��c���   ���   �Ѓ�;�����_^[���   ;�������]���������������������������U����   SVW��@����0   ������E�8 t ��E�Q��c�B�H�у�;��*����E�     _^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ��c�B��  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   ������} t�E�x��u�   �3�_^[��]��������������������U����   SVW��4����3   ������}s�E   �E��P������E��}� u3��:�} t�E��Pj �M�Q������E�� �����E����E���c   �E�_^[���   ;�������]��������������������������������������������U����   SVW��<����1   ������=�c tE�}sǅ<���   �	�E��<�����j j ��<���Q��c�B��H  �у�;������j�EP������_^[���   ;��������]���������������������������������������������������U����   SVW��<����1   ������=�c tE�}sǅ<���   �	�E��<�����j j ��<���Q��c�B��H  �у�;��F����j�EP�+����_^[���   ;��&�����]���������������������������������������������������U����   SVW��<����1   ������=�c tE�}sǅ<���   �	�E��<�����j j ��<���Q��c�B��H  �у�;������j�EP�k����_^[���   ;��f�����]���������������������������������������������������U����   SVW��<����1   ������=�c tI�}sǅ<���   �	�E��<�����MQ�UR��<���P��c�Q��H  �Ѓ�;�������j�EP�����_^[���   ;�������]�����������������������������������������������U����   SVW��<����1   ������=�c ��   �} tK�}sǅ<���   �	�E��<�����MQ�UR��<���P��c�Q��H  �Ѓ�;�������[�I�}sǅ<���   �	�E��<�����MQ�UR��<���P��c�Q���  �Ѓ�;�������EP�MQ�����_^[���   ;�������]������������������������������������������������������������������������U����   SVW��<����1   ������=�c tE�}sǅ<���   �	�E��<�����j j ��<���Q��c�B��H  �у�;�������j�EP� ����_^[���   ;�������]���������������������������������������������������U����   SVW��<����1   ������=�c tI�}sǅ<���   �	�E��<�����MQ�UR��<���P��c�Q��H  �Ѓ�;������j�EP�������_^[���   ;��������]�����������������������������������������������U����   SVW��<����1   ������=�c ��   �} tK�}sǅ<���   �	�E��<�����MQ�UR��<���P��c�Q��H  �Ѓ�;��H����[�I�}sǅ<���   �	�E��<�����MQ�UR��<���P��c�Q���  �Ѓ�;��������EP�MQ�������_^[���   ;��������]������������������������������������������������������������������������U����   SVW��4����3   ������} tG�E�E��=�c t�E�x��u�E��P�\��������E�P��c�Q�B�Ѓ�;��%���_^[���   ;�������]����������������������������������U����   SVW��4����3   ������} tG�E�E��=�c t�E�x��u�E��P���������E�P��c�Q�B�Ѓ�;�����_^[���   ;��u�����]����������������������������������U����   SVW��@����0   ������EP�������_^[���   ;�������]�������������������U����   SVW��@����0   ������EP������_^[���   ;��������]�������������������U����   SVW��4����3   ������E��8�����8���Q������_^[���   ;��j�����]�����������������������U����   SVW��4����3   ������E��8�����8���Q������_^[���   ;��
�����]�����������������������U����   SVW��4����3   ������E��8�����8���Q������_^[���   ;�������]�����������������������U����   SVW��4����3   ������E��8�����8���Q�t����_^[���   ;��J�����]�����������������������U����   SVW��@����0   �������EP��c�Q|��Ѓ�;������_^[���   ;��������]����������������������������������U����   SVW��@����0   �������h   ��c�H|��҃�;�����_^[���   ;��u�����]����������������������������������U����   SVW��@����0   ������E�8 t ��E�Q��c�B|�H�у�;��
����E�     _^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H|�Q�҃�;�����_^[���   ;��x�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H|�Q�҃�;�����_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H|�Q�҃�;�����_^[���   ;��x�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B|�H�у�;�����_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVW��@����0   ������E�M�H4�E�@���E�@8���E�@<���E�@@��E�@D���E�@H���E�@L9��E�@P���E�@h��E�@pg��E�@X~��E�@\Ͽ�E�@`o��E�@d���E�@Tʿ�E�@l���E�M�H �E�M��E�M�H0�E�M�H(�E�@,    _^[��]����������������������������������������������������������������������U���h  SVW�������Z   ������j h�   ��\���P�H�����j �EP�MQ�UR�EP��\���Q��������E �E�h�   ��\���P�MQ�URj�b����R��P��	����XZ_^[��h  ;��6�����]Ë�   ��	\����   �	np ��������������������������������������������������������̋�`<����������̋�`����������̋�` ����������̋�`0����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`����������̋�`����������̋�`,�����������U����   SVW��@����0   �����󫡨c�HL��8  ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;��R����E�     _^[���   ;��9�����]��������������������������������������U����   SVW��@����0   �����󫡨c�HL����;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;��r����E�     _^[���   ;��Y�����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL���   �Ѓ�;������_^[���   ;��������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HL���   �҃�;��u���_^[���   ;��e�����]� �������������������������������U����   SVW��@����0   �����󫡨c�HL��Q��;�����_^[���   ;��������]�������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;������E�     _^[���   ;�������]��������������������������������������U����   SVWQ������;   ������Y�XD3ŉE��M�M��������E�P�MQ�U�R��c�HL�Q�҃�;������E�P�M����M��H����ER��P�d�	�Q���XZ_^[�M�3��>������   ;��������]� ��   l�	����   x�	bc �����������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BL��   �у�;��(���_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HL�Q�҃�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL�B �Ѓ�;��/���_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL�B$�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL�B(�Ѓ�;��O���_^[���   ;��?�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HL�Q,�҃�;������_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�QL�B0�Ѓ�;��S���_^[���   ;��C�����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��c�BL�H4�у�;������_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL�B8�Ѓ�;��_���_^[���   ;��O�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL�B<�Ѓ�;������_^[���   ;��������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL���   �Ѓ�;��|���_^[���   ;��l�����]�������������������������U����   SVWQ������:   ������Y�M���E�P�����Q��c�BL��   �у�;�����P�M���������G����E_^[���   ;��������]� ����������������������������������������U����   SVWQ������:   ������Y�M���EP�M�Q�����R��c�HL��T  �҃�;��b���P�M��������������E_^[���   ;��;�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL�B@�Ѓ�;������_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���j �E�P��c�QL�BD�Ѓ�;��]���_^[���   ;��M�����]��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��c�BL�M����   ��;������_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��c�BL�M����   ��;��h���_^[���   ;��X�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��c�BL�M���4  ��;������_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��c�BL�M����   ��;��h���_^[���   ;��X�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��c�BL�M����   ��;������_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��c�BL�M���  ��;��h���_^[���   ;��X�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP��c�QL�M����   ��;������_^[���   ;��������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��c�QL�M����   ��;��|���_^[���   ;��l�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��c�QL�M���0  ��;�����_^[���   ;��������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BL�HT�у�;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HL�QX�҃�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���j �EP�M�Q��c�BL�H\�у�;��)���_^[���   ;�������]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j �EP�M�Q��c�BL�H`�у�;�����_^[���   ;�������]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j�EP�M�Q��c�BL�H\�у�;��)���_^[���   ;�������]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j�EP�M�Q��c�BL�H`�у�;�����_^[���   ;�������]� �����������������������������������U���$  SVWQ�������I   ������Y�M��M������h�  �������3���P����������j �E�P������Q�M��R���������������������(�����������tǅ���    �M��;����������M������������M����������R��P���	����XZ_^[��$  ;�������]Ë�   ��	����   ��	dat ����������������������������������������������������������������������������U���   SVWQ�� ����@   ������Y�M�j���������h�  ��$��������P������;���j�����P�����Q�M������������������������_^[��   ;�������]���������������������������������������������������U���   SVWQ�� ����@   ������Y�M��EP���������h�  ��$����,���P������y���j�����Q�����R�M������������+���������P���_^[��   ;��������]� ����������������������������������������������U���   SVWQ�� ����@   ������Y�M��EP������]���h�  ��$����l���P���������j�����Q�����R�M��3���������k������������_^[��   ;��$�����]� ����������������������������������������������U���  SVWQ�������C   ������Y�M��M��~���h�  ���������P������ ���j �E�P�����Q�M����������������������������������t�M������M������E��M�����P�M������M������ER��P��	袾��XZ_^[��  ;�������]� �   �	����   �	dat ����������������������������������������������������������������U���  SVWQ�������C   ������Y�M��M��N���h�  ���������P����������j �E�P�����Q�M����������������������x�����������t�M������M������E��M������P�M�����M��o����ER��P�8�	�r���XZ_^[��  ;��������]� �   @�	����   L�	dat ����������������������������������������������������������������U���$  SVWQ�������I   ������Y�M��M�����h�  �������S���P����������j �E�P������Q�M��r���������������������H�����������t��ٝ����M��]���م�����M��~���ٝ����M��?���م���R��P�h�	�?���XZ_^[��$  ;�������]�   p�	����   |�	dat ����������������������������������������������������������������U���$  SVWQ�������I   ������Y�M��M�����h�  �������#���P�������p���j �E�P������Q�M��B��������������������������������tǅ���    �M��+����������M�����������M����������R��P���	����XZ_^[��$  ;�������]Ë�   ��	����   ��	dat ����������������������������������������������������������������������������U���  SVWQ�������C   ������Y�M��M�讳��h�  ����������P������0���j �E�P�����Q�M����������������������������������t�M�����M�������E� �M��������P�E��P�M�������ER��P���	�ι��XZ_^[��  ;��K�����]� �   ��	����   ��	dat ����������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E�����E����X�E�_^[��]���������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL��  �Ѓ�;��L���_^[���   ;��<�����]�������������������������U����   SVWQ��$����7   ������Y�M���j�EP�M�Q��(���R��c�HL��  �҃�;��������P�E��P�E_^[���   ;�������]� ������������������������������������������U����   SVWQ��$����7   ������Y�M���j �EP�M�Q��(���R��c�HL��  �҃�;��0�����P�E��P�E_^[���   ;�������]� ������������������������������������������U���  SVWQ�������C   ������Y�M��M��n���h�  ���������P����������j �E�P�����Q�M����������������������������������t�M�f����M������E� �M�������P�E��P�M������ER��P��	莶��XZ_^[��  ;�������]� �   $�	����   0�	dat ����������������������������������������������������������������������������U���  SVWQ�������C   ������Y�M��M��.���h�  ������c���P���������j �E�P�����Q�M����������������������X�����������t�M�&����M��m����E� �M��r�����P�E��P�M��K����ER��P�\�	�N���XZ_^[��  ;��������]� �   d�	����   p�	dat ����������������������������������������������������������������������������U���  SVWQ�������C   ������Y�M��M�����h�  ������#���P������p���j �E�P�����Q�M��B�������������������������������t�M������M��-����E� �M��2�����P�E��P�M������ER��P���	����XZ_^[��  ;�������]� �   ��	����   ��	dat ����������������������������������������������������������������������������U���$  SVWQ�������I   ������Y�M��M�讬��h�  �����������P�������0���j �E�P������Q�M�����������������������������������tǅ���    �M�������������M��q���������M�����������R��P���	�Ͳ��XZ_^[��$  ;��J�����]Ë�   ��	����   ��	dat ����������������������������������������������������������������������������U���   SVWQ�� ����@   ������Y�M�Q�E�$���������h�  ��$�������P����������j�����P�����Q�M��`���������������������_^[��   ;��Q�����]� �������������������������������������������U���   SVWQ�� ����@   ������Y�M��EP����������h�  ��$��������P������)���j�����Q�����R�M��������������������� ���_^[��   ;�蔽����]� ����������������������������������������������U���   SVWQ�� ����@   ������Y�M��EP������1���h�  ��$�������P������i���j�����Q�����R�M���������������������@���_^[��   ;��Լ����]� ����������������������������������������������U���   SVWQ�� ����@   ������Y�M��EP������q���h�  ��$����\���P���������j�����Q�����R�M��#���������[������������_^[��   ;�������]� ����������������������������������������������U���   SVWQ�� ����@   ������Y�M��EP���������h�  ��$�������P����������j�����Q�����R�M��c����������������������_^[��   ;��T�����]� ����������������������������������������������U���   SVWQ�� ����@   ������Y�M��EP����������h�  ��$��������P������)���j�����Q�����R�M��������������������� ���_^[��   ;�蔺����]� ����������������������������������������������U���   SVWQ�� ����@   ������Y�M��EP����������h�  ��$�������P������i���j�����Q�����R�M���������������������@���_^[��   ;��Թ����]� ����������������������������������������������U���  SVWQ�������C   ������Y�M��M��.���h�  ������c���P���������j �E�P�����Q�M����������������������X�����������t�M�&����M��m����E� �M��r�����P�E��P�M��K����ER��P�\�	�N���XZ_^[��  ;��˸����]� �   d�	����   p�	dat ����������������������������������������������������������������������������U���$  SVWQ�������I   ������Y�M��M�����h�  �������#���P�������p���j �E�P������Q�M��B��������������������������������tǅ���    �M��+����������M�����������M����������R��P���	����XZ_^[��$  ;�芷����]Ë�   ��	����   ��	dat ����������������������������������������������������������������������������U���$  SVWQ�������I   ������Y�M��M�讣��h�  �����������P�������0���j �E�P������Q�M�����������������������������������tǅ���    �M�������������M��q���������M�����������R��P���	�ͩ��XZ_^[��$  ;��J�����]Ë�   ��	����   ��	dat ����������������������������������������������������������������������������U����   SVWQ��$����7   ������Y�M��M�������E�}�t�}�t�}�tǅ$���    �
ǅ$���   ��$���_^[���   ;��t�����]���������������������������������U���   SVWQ�� ����@   ������Y�M��EP������!���h�  ���������P��(����Y���j�����Q��(���R�M��������(�������������0���_^[��   ;��Ĵ����]� ����������������������������������������������U���   SVWQ�� ����@   ������Y�M��EP������A���h�  ��$����L���P���������j�����Q�����R�M�����������K���������p���_^[��   ;�������]� ����������������������������������������������U���   SVWQ�� ����@   ������Y�M��EP���������h�  ��$�������P����������j�����Q�����R�M��S���������������������_^[��   ;��D�����]� ����������������������������������������������U����   SVW��@����0   �������EP��c�Q���   �Ѓ�;��Ѳ��_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP��c�Q���   �Ѓ�;��a���_^[���   ;��Q�����]������������������������������U����   SVW��@����0   �����󫡨c�H���   ��;������_^[���   ;�������]����������������������U����   SVW��@����0   �����󫡨c�H���   ��;�虱��_^[���   ;�艱����]����������������������U����   SVW��@����0   �������E�Q��c�B���   �у�;��/����E�     _^[���   ;�������]�����������������������������������U����   SVW��@����0   �������EP��c�Q���   �Ѓ�;�豰��_^[���   ;�衰����]������������������������������U����   SVW��4����3   �����������E��}� u3��_��EP�MQ�UR�E�P��c�Q��@  �Ѓ�;��#�����u+�}� t��E�P��c�Q@�BH�Ѓ�;�������E�    �E�_^[���   ;�������]����������������������������������������������U����   SVW��@����0   �������EP�M�� Q�UR�EP��c�Q��@  �Ѓ�;��b���_^[���   ;��R�����]�������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��c�Q���   �Ѓ�;�����_^[���   ;��ծ����]����������������������������������U����   SVW��@����0   �������E0P�M,Q�U(R�E$P�M Qj �UR�EP�MQ�UR�EP�MQ��c�B���   �у�0;��G���_^[���   ;��7�����]������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL�Bd�Ѓ�;��ϭ��_^[���   ;�迭����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL�Bh�Ѓ�;��_���_^[���   ;��O�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HL�Ql�҃�;�����_^[���   ;��ج����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BL��  �у�;��h���_^[���   ;��X�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL�Bt�Ѓ�;�����_^[���   ;��߫����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�QL���   �Ѓ�;��p���_^[���   ;��`�����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�QL�B|�Ѓ�;�����_^[���   ;�������]� �����������������������������U���`  SVWQ�������X   ������Y�XD3ŉE��M������E�}� u3��  �E�    �E�    �E�    �M��$�����|����n����E艅|����E��E��EPh]  �M�����j j �E�P�M�������u��   �M��z����E���E܉Eă}� ��   �M������E܋EĉE���|���Ph�   �ל������u�   �}� u�   j �M������EЃ}� u�l�E�P�M��2����E�P�/������}� t��E�P��c�Q@�BH�Ѓ�;��v����E�    �Z����E艅������|��������M�褙���������Z�}� t��E�P��c�Q@�BH�Ѓ�;��"����E�    �E�P褭����ǅ����    ��|���������M��H���������R��P�h�	�N���XZ_^[�M�3��;�����`  ;��������]� �I    p�	����   ��	|���$   ��	cd ctr �������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E��@    �E��@    �E��@     �E��@   �E��@    �E�_^[��]�������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��c���   �M��B��;�����_^[���   ;��������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP��c���   �M����   ��;�艦��_^[���   ;��y�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP��c���   �M��B<��;�����_^[���   ;��������]� ����������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL���   �Ѓ�;�蜥��_^[���   ;�茥����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL���   �Ѓ�;��,���_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BL���   �у�;�踤��_^[���   ;�訤����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL���   �Ѓ�;��<���_^[���   ;��,�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BL���   �у�;��ȣ��_^[���   ;�踣����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BL���   �у�;��H���_^[���   ;��8�����]� ����������������������������������U����   SVW��@����0   ������E���M���;��ݢ��_^[���   ;��͢����]��������������������������U����   SVW��@����0   �������EP�M��M�B��;��x���_^[���   ;��h�����]���������������������U����   SVW��@����0   �������EP�MQ�U��M�P��;�����_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�M��M�B��;�蜡��_^[���   ;�茡����]�������������������������U����   SVWQ��4����3   ������Y�M��E��M�H�E��M�H��hI�h��h�h���E��HQ�UR�EPQ�E�$�MQ�U��BP�M�Q��c�BL���   �у�,;�����_^[���   ;��ՠ����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL���   �Ѓ�;��\���_^[���   ;��L�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BL���   �у�;�����_^[���   ;��؟����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BL���   �у�;��h���_^[���   ;��X�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BL���   �у�;�����_^[���   ;��؞����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BL���   �у�;��h���_^[���   ;��X�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BL���   �у�;�����_^[���   ;��؝����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QL��<  �Ѓ�;��l���_^[���   ;��\�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R��c�HL��@  �҃�;�����_^[���   ;��ٜ����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�QL��D  �Ѓ�;��`���_^[���   ;��P�����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��c�BL��H  �у�;��ܛ��_^[���   ;��̛����]� ��������������������������������������U���  SVW�������D   ������M�蒵���M��y����} t�M�辴����u"ǅ����   �M��Q����M������������Qj�M�莴��P�M������M��}����E�E�E؍E�Ph=���������� ����M�������M�蹢���� ���R��P�X�	�O���XZ_^[��  ;��̚����]�   `�	����$   �	����   x�	active mu ������������������������������������������������������������������������������U���  SVW�������D   ������M��B����M��)����} t�M��n�����u"ǅ����   �M������M�輡���������Qj�M��>���P�M�|����M��-����E�E�E؍E�Ph<��赌������ ����M�讂���M��i����� ���R��P���	�����XZ_^[��  ;��|�����]�   ��	����$   ��	����   ��	active mu ������������������������������������������������������������������������������U����   SVW��@����0   �������EP�MQ�UR��c�HL��$  �҃�;�躘��_^[���   ;�誘����]�����������������������U����   SVW��@����0   �������EP�MQ��c�BL��(  �у�;��M���_^[���   ;��=�����]��������������������������U����   SVW��@����0   �������EP�MQ��c�BL��,  �у�;��ݗ��_^[���   ;��͗����]��������������������������U����   SVW��@����0   �����󫡨c�HL��\  ��;��y���_^[���   ;��i�����]����������������������U����   SVWQ��4����3   ������Y�M�艳���M���E�_^[���   ;�������]�����������������������������U����   SVW��@����0   �����󫡨c���   �􋑌   ��;�趖��_^[���   ;�視����]�����������������������������������U����   SVWQ��4����3   ������Y�M��E�P�������E��     _^[���   ;��8�����]���������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E�M��;t3��M�E�x t�E��x t�E�M��P;Qt3��)�E�x t�E��x t�E�M��P;Qt3���   _^[��]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M����������_^[���   ;�������]� ��������������������U����   SVWQ��(����6   ������Y�M��E�    �	�E���E�E�P�M��&����8 t��E�_^[���   ;��u�����]����������������������������������U����   SVWQ��$����7   ������Y�M��E�    �	�E���E�E�P�M�覓���8 t$�E�P�M�蕓�����M�Q�M臓���;t��} t�E�M��}� ~�E�P�M��]����8 uǅ$���   �
ǅ$���    ��$���_^[���   ;�蕓����]� ���������������������������������������������������������������U����   SVW��4����3   ������j�k   ���E��}� t	�E��x u3�� ��EP�MQ�UR�E��H�у�;�����_^[���   ;�������]�������������������������������U����   SVW��@����0   ������h�c�EPhD ������_^[���   ;��|�����]�������������������������U����   SVWQ��(����6   ������Y�M�j\�v������E�}� t	�E�x\ u���E�P�M�Q\�҃�;������E�_^[���   ;��������]���������������������������������U����   SVWQ��(����6   ������Y�M�j\��������E�}� t	�E�x\ u�$��E�P�M�Q\�҃�;��w����EP�M������E�_^[���   ;��X�����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�j\�F������E�}� t	�E�x\ u�$��E�P�M�Q\�҃�;��א���EP�M������E�_^[���   ;�踐����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�j\�������E�}� t	�E�x\ u�0��E�P�M�Q\�҃�;��7����EP�M��p����EP�M��,����E�_^[���   ;�������]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�j\��������E�}� t	�E�x\ u�<��E�P�M�Q\�҃�;�臏���EP�M�������EP�M��|����EP�M��p����E�_^[���   ;��P�����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�j`�6������E�}� t	�E�x` u���E�P�M�Q`�҃�;��ǎ��_^[���   ;�跎����]������������������������������������U����   SVWQ��(����6   ������Y�M�jd�������E�}� t	�E�xd u���EP�M�Q�U�Bd�Ѓ�;��3���_^[���   ;��#�����]� �����������������������������U����   SVWQ��(����6   ������Y�M�jh�������E�}� t	�E�xh u���EP�M�Q�U�Bh�Ѓ�;�裍��_^[���   ;�蓍����]� �����������������������������U����   SVWQ��(����6   ������Y�M�jl�������E�}� t	�E�xl u���E�P�M�Ql�҃�;�����_^[���   ;�������]������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;��x���_^[���   ;��h�����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h�   �S������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;��؋��_^[���   ;��ȋ����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�jp�������E�}� t	�E�xp u��c���EP�M�Q�U�Bp�Ѓ�;��>���_^[���   ;��.�����]� ����������������������������������������U����   SVWQ������:   ������Y�M�jt�������E�}� t	�E�xt uh�c�M�����E�:��EP�M�Q�����R�E�Ht�у�;�茊��P�M�W��������褳���E_^[���   ;��e�����]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�jx�F������E�}� t	�E�xx u�E����E�P�MQ�U�Bx�Ѓ�;��Љ���E�_^[���   ;�轉����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�jx�������E�}� t	�E�x| u3����E�P�MQ�U�B|�Ѓ�;��1���_^[���   ;��!�����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jx�������E�}� t	�E�x| u�   �#��E�P�MQ�U�B|�Ѓ�;�莈�������_^[���   ;��w�����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVW��4����3   ������j�+������E��}� t	�E��x u3���E���H��;������_^[���   ;�豇����]������������������������������U����   SVW��4����3   ������E�8 u�?j�������E��}� t	�E��x u�!��EP�M��Q�҃�;��2����E�     _^[���   ;�������]��������������������������������������U����   SVWQ��(����6   ������Y�M��} u3��@j��������E�}� t	�E�x u3�� ��EP�MQ�U�R�E�H�у�;�胆��_^[���   ;��s�����]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M�j�V������E�}� t	�E�x u3����EP�M�Q�U�B�Ѓ�;�����_^[���   ;��х����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3����EP�M�Q�U�B�Ѓ�;��A���_^[���   ;��1�����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j �������E�}� t	�E�x  u3����E�P�M�Q �҃�;�襄��_^[���   ;�蕄����]����������������������������������U����   SVWQ��(����6   ������Y�M�j$�������E�}� t	�E�x$ u3����E�P�M�Q$�҃�;�����_^[���   ;�������]����������������������������������U����   SVWQ��(����6   ������Y�M�j(��������E�}� t	�E�x( u3��$��EP�MQ�UR�E�P�M�Q(�҃�;��y���_^[���   ;��i�����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j,�V������E�}� t	�E�x, u3�� ��EP�MQ�U�R�E�H,�у�;��݂��_^[���   ;��͂����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�j(�������E�}� t	�E�x0 u3��$��EP�MQ�UR�E�P�M�Q0�҃�;��9���_^[���   ;��)�����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j4�������E�}� t	�E�x4 u3����E�P�M�Q4�҃�;�襁��_^[���   ;�蕁����]����������������������������������U����   SVWQ��(����6   ������Y�M�j8�������E�}� t	�E�x8 u3��(��EP�MQ�UR�EP�M�Q�U�B8�Ѓ�;�����_^[���   ;��������]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�j<��������E�}� t	�E�x< u���EP�M�Q�U�B<�Ѓ�;��c���_^[���   ;��S�����]� �����������������������������U����   SVWQ��(����6   ������Y�M�jD�F������E�}� t	�E�xD u3����E�P�M�QD�҃�;�����_^[���   ;�������]����������������������������������U����   SVWQ��(����6   ������Y�M�jH�������E�}� u���EP�M�Q�U�BH�Ѓ�;��L��_^[���   ;��<����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�jL�&������E�}� u3����EP�M�Q�U�BL�Ѓ�;��~��_^[���   ;��~����]� ������������������������������������U����   SVWQ��(����6   ������Y�M�jP�������E�}� u3�� ��EP�MQ�U�R�E�HP�у�;��&~��_^[���   ;��~����]� ��������������������������������U����   SVWQ��(����6   ������Y�M�jT�������E�}� u3����E�P�M�QT�҃�;��}��_^[���   ;��}����]���������������������������U����   SVWQ��(����6   ������Y�M�jX�������E�}� u���EP�M�Q�U�BX�Ѓ�;��}��_^[���   ;��}����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� u3��/��EP�MQ�UR�EP�MQ�U�R�E싈�   �у�;��t|��_^[���   ;��d|����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �C������E�}� u3��'��EP�MQ�UR�E�P�M싑�   �҃�;���{��_^[���   ;��{����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� u3����EP�M�Q�U싂�   �Ѓ�;��4{��_^[���   ;��${����]� ������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� u3����EP�M�Q�U싂�   �Ѓ�;��z��_^[���   ;��z����]� ������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� u3����EP�M�Q�U싂�   �Ѓ�;��z��_^[���   ;��z����]� ������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� u�'��EP�MQ�UR�E�P�M싑�   �҃�;��~y��_^[���   ;��ny����]� ����������������������������������������U����   SVW������9   ������h�   �X������E��}� u�M�B����E�9��EP�� ���Q�U����   �Ѓ�;���x��P�M�օ���� ����8����E_^[���   ;��x����]���������������������������������������������������U����   SVWQ������?   ������Y�M�h�   �������E�}� t�E샸�    uj ������,���P�M�|����E�9��EP�����Q�U�M����   ��;���w��P�M�ɔ������������E_^[���   ;���w����]� �������������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;��4w��_^[���   ;��$w����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����EP�U�M����   ��;��v��_^[���   ;��|v����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� t�E샸�    u3����EP�U�M����   ��;���u��_^[���   ;���u����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3����EP�U�M����   ��;��Lu��_^[���   ;��<u����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �#������E�}� t�E샸�    u3����E�M����   ��;��t��_^[���   ;��t����]���������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;��t��_^[���   ;���s����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u���EP�U�M����   ��;��^s��_^[���   ;��Ns����]� ����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �3������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;��r��_^[���   ;��r����]� ����������������������������������������������U����   SVW������;   ������XD3ŉE��EP�M��J����EP�4v�����E؃}� t��E�P�U؋E؋H �RL��;��r���E�P�M萛���M��Nb���ER��P�\%
�We��XZ_^[�M�3��D������   ;���q����]Ë�   d%
����   p%
bc �������������������������������������������������������������U���  SVWQ�������A   ������Y�XD3ŉE��M�j h�  �M��Xu���} u�   �oj h�  �M��7k���E�}� u3��S�M���]���EPh�  �M��j��Q�E�$h�  �M���^��j �E�P�M��j��ǅ ���   �M��a���� ���R��P��&
�d��XZ_^[�M�3�������  ;��p����]� �I    �&
����   �&
bc �����������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H@�Qd�҃�;���o��_^[���   ;���o����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$�E�P��c�QH�B �Ѓ�;��Xo��_^[���   ;��Ho����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH���   �у�;���n��_^[���   ;���n����]� ����������������������������������U���  SVWQ�������A   ������Y�M���E�P�� ���Q��c�BH�HP�у�;��Xn���   ���}�E_^[��  ;��9n����]� �����������������������������������U���  SVWQ�������A   ������Y�M���E�P�� ���Q��c�BH�HT�у�;���m���   ���}�E_^[��  ;��m����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH���  �у�;��8m��_^[���   ;��(m����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH��   �у�;��l��_^[���   ;��l����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HH��D  �҃�;��5l��_^[���   ;��%l����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HH��H  �҃�;��k��_^[���   ;��k����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH���  �Ѓ�;��<k��_^[���   ;��,k����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH���  �у�;���j��_^[���   ;��j����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���j �E�P��c�QH�Bd�Ѓ�;��Mj��_^[���   ;��=j����]��������������������������U����   SVWQ��4����3   ������Y�M���EPj �M�Q��c�BH�Hh�у�;���i��_^[���   ;���i����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j�E�P��c�QH�Bd�Ѓ�;��]i��_^[���   ;��Mi����]��������������������������U����   SVWQ��4����3   ������Y�M���EPj�M�Q��c�BH�Hh�у�;���h��_^[���   ;���h����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j�E�P��c�QH�Bd�Ѓ�;��mh�������_^[���   ;��Wh����]������������������������������������U����   SVWQ��4����3   ������Y�M���EPj�M�Q��c�BH�Hh�у�;���g��_^[���   ;���g����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HH���   �҃�;��eg��_^[���   ;��Ug����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HH���   �҃�;���f��_^[���   ;���f����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH�Bt�Ѓ�;��of��_^[���   ;��_f����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R��c�HH���  �҃�;���e��_^[���   ;���e����]� �����������������������������������U����   SVWQ��(����6   ������Y�M��EP�u�����E�}� t�EP�M�Q�M��BT���E�_^[���   ;��Ue����]� �������������������������������U����   SVWQ��(����6   ������Y�M��EP�MQ��w�����E�}� t�EP�M�Q�M��S���E�_^[���   ;���d����]� ���������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��  �Ѓ�;��ld��_^[���   ;��\d����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��  �Ѓ�;���c��_^[���   ;���c����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH��  �у�;��c��_^[���   ;��xc����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH��  �у�;��c��_^[���   ;���b����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HH��P  �҃�;��b��_^[���   ;��ub����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HH��  �҃�;��b��_^[���   ;���a����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH���  �Ѓ�;��a��_^[���   ;��|a����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH���  �Ѓ�;��a��_^[���   ;��a����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH���  �Ѓ�;��`��_^[���   ;��`����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��   �Ѓ�;��<`��_^[���   ;��,`����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��$  �Ѓ�;���_��_^[���   ;��_����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HH��(  �҃�;��U_��_^[���   ;��E_����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�QH��,  �Ѓ�;���^��_^[���   ;���^����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH��<  �у�;��X^��_^[���   ;��H^����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��t  �Ѓ�;���]��_^[���   ;���]����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HH��@  �҃�;��e]��_^[���   ;��U]����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH��h  �у�;���\��_^[���   ;���\����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�j h�  �M�� y�����l����E�M���v�����}�u�E���3�_^[���   ;��H\����]�������������������������������������U����   SVWQ��4����3   ������Y�M�j h�  �M��x�����mX��_^[���   ;���[����]��������������������U����   SVWQ�� ����8   ������Y�M���EP�MQQ�E�$�U�R��$���P��c�QH��,  �Ѓ�;��f[���M���P�Q�@�A�E_^[���   ;��@[����]� ������������������������������������������U����   SVWQ�� ����8   ������Y�M���EP�MQQ�E�$�U�R��$���P��c�QH��0  �Ѓ�;��Z���M���P�Q�@�A�E_^[���   ;��Z����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HH��4  �҃�;��Z��_^[���   ;��Z����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��8  �Ѓ�;��Y��_^[���   ;��Y����]�������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$�E�P��c�QH��<  �Ѓ�;��%Y��_^[���   ;��Y����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��@  �Ѓ�;��X��_^[���   ;��X����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HH��D  �҃�;��5X��_^[���   ;��%X����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EPQ�E�$�MQ�U�R��c�HH��H  �҃�;��W��_^[���   ;��W����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH���  �Ѓ�;��,W��_^[���   ;��W����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��L  �Ѓ�;��V��_^[���   ;��V����]�������������������������U����   SVWQ��4����3   ������Y�M��E��     �E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M���j�E��Q��c�BH���  �у�;���U��_^[���   ;���U����]�������������������������������������U����   SVWQ��4����3   ������Y�M���EP��c�QH���  �Ѓ�;��|U���M���E�3Ƀ8 ����_^[���   ;��ZU����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���j �E��Q��c�BH���  �у�;���T��_^[���   ;���T����]�������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��h  �Ѓ�;��lT��_^[���   ;��\T����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��l  �Ѓ�;���S��_^[���   ;���S����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��p  �Ѓ�;��S��_^[���   ;��|S����]�������������������������U����   SVWQ�� ����8   ������Y�M���E�P��$���Q��c�BH��t  �у�;��S���U��
�H�J�@�B�E_^[���   ;���R����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��x  �Ѓ�;��|R��_^[���   ;��lR����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH��|  �у�;��R��_^[���   ;���Q����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$�E�P��c�QH���  �Ѓ�;��Q��_^[���   ;��uQ����]� �������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$�E�P��c�QH���  �Ѓ�;��Q��_^[���   ;���P����]� �������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$�E�P��c�QH���  �Ѓ�;��P��_^[���   ;��uP����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH���  �у�;��P��_^[���   ;���O����]� ����������������������������������U����   SVW��@����0   �������EP�MQQ�E�$�UR�EP�MQ��c�BH���   �у�;��zO��_^[���   ;��jO����]���������������������������������������U����   SVW��@����0   �������EPQ�E�$�MQ�UR�EP��c�QH���   �Ѓ�;���N��_^[���   ;���N����]���������������������������U����   SVW��@����0   �������E�M�8O�p���E�EP�MQ�UR�F]����_^[���   ;��jN����]�����������������������U����   SVW��@����0   ������E;E}�E��E;E~�E��E_^[��]�������������������������������U���,  SVW��������   ������M�#h���E��E�    �M��o���E��E�    �E�    �E�    �E�    �}� u
�   ��  �M��V��=�  ��	  j h:  �M��N���E��M�HC���E�ǅP���    �M�S����,����M�e:���� ����M�L�������������j���E�    �	�E����E��E�;E���   �� ��� ��   j��E�P�� �����U����t�����t����tk��t���k������HQ��9E�t룋�t���k������M��������������;�P���~��������P�����t���k������?��EԉE��6�E����M�����,�����,����D;Du�Eԃ��E��	�Eԃ��E������}� tj �EP�M��@����u
�2  �-  �}� tz�M���W����tn�M��A��;E�ua��hT�hB��%P�M�k�Q��c�B��H  �у�;��K���E��}� u
��  ��  �E�k�P�M�Q�M��WW��P�N������hT�hB��)P�M�k�Q��c�B��H  �у�;��UK���E��}� u
�m  �h  �E�k�P�M�Q�U�R�M������P��� ~K��hT�hB��.P��P�������Q��c�B��H  �у�;���J���E��}� u
�  ��
  j��E�P�M�wG����u
��
  ��
  �}� tj�EP�M��??����u
��
  �
  �}� t�M��Qa���������
ǅ����    �������E��M�l���E��E�    �E�    �	�E����E��E�;E��/  �� ��� ��  j��E�P�� ����(S����t�����t������  ��t���k������N��9E�t�ǅ\���    ǅh���    ���h�������h�����t���k������VT��9�h�����  ��h���P��t���k������M����u밋�h���P��t���k������r6����D�����D�������\����U���,��������\�������\�����D�������\����U�����\�������\�����D�������\����U���,����D����\�������\�����D�����   ��\����E�����\�������\�����D�������\����U���,����D����\�������\�����D�����   ��\����E�����\�������\�����D�������\����U���,����D����\�������\�����D�����   ��\����E�����\�������\����7�����\��������������� ��  j�������+���P�E�P������?3��ǅ\���    ��\����M����������}� t%������k�E��M�k�M����P�Q�@�A������k�E��M�k�Mȋ��P�Q�@�A��\���;�������   ��\����M���;�������   ��\����M��D���������D�����\����M��T�����8�����8���������������wj�������$�X
��D�������,����Uԉ�F��D�������,����UԉT�.��D�������,����UԉT���D�������,����UԉT��\�������\��������Eԃ��Eԋ�\���;�����������N  �E����M�����,�����,����D3�;D�U��}� ��   �E�����,����k�U��E�k�E��
��J�H�R�P�E�����,����Tk�U��Eԃ�k�E��
��J�H�R�P�E�����,����Tk�U��Eԃ�k�E��
��J�H�R�P�}� t2�E�����,����Tk�U��Eԃ�k�E��
��J�H�R�P�E�����,����k�U��E�k�Eȋ
��J�H�R�P�E�����,����Uԉ�Eԃ��EԋE�����,����Tk�U��E�k�Eȋ
��J�H�R�P�E�����,����UԉT�Eԃ��EԋE�����,����Tk�U��E�k�Eȋ
��J�H�R�P�E�����,����UԉT�Eԃ��Eԃ}� tM�E�����,����Tk�U��E�k�Eȋ
��J�H�R�P�E�����,����UԉT�Eԃ��E�� �E����M�����,�����,����D�D
�����E�P�w>�����E�P�k>�����  �M�=M��=  ��  �M�>\���������M��Y���������E�    �	�E����E��E�;�����}?�E��������|� t�E����������EԍP�M���E����������EԍLP��M�뭋�hT�hB�   P�M�k�Q��c�B��H  �у�;��5C���E��}� u3��q  �E�k�P�M�Q�U�R�E������hT�hB�   P��������Q��c�B��H  �у�;���B�������������� u3��  ��������P������Q������R�.E�����Eԙ+���P�E�P�M��Z����u"�E�P��<����������P��<����3��  �M�d���EȋM�Z��������ǅ����    ǅ����    �E�    �	�E����E��E�;�������  ǅ����    ������������������������M�������;���   ��������;E�}�������������T;U�|hT�hB�   P�y1�����   �����������k�E�������k�Mȋ��P�Q�@�A���������������������������Tk�U�������k�Eȋ
��J�H�R�P�������������������E��������|� ��   ��������;E�}�����������;E�|hT�hB�   P�0�����   �����������k�E�������k�Mȋ��P�Q�@�A��������������������k�E�������k�Mȋ��P�Q�@�A���������������E�������������������������E�    �	�E����E��Eԙ+���9E�}#�E��������D�    �E���������   �Ǎ�����P�_:�����E�P�S:�����   �&�E�P�@:�����E�P�4:�����E�P�(:����3�R��P��W
�3��XZ_^[��,  ;��?����]ÍI    �W
����   �W
����   �W
����   �W
���   �W
����   �W
osadr pointsort ngonpointmap opadr sttpadr �+P
BP
ZP
rP
��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������} t �} t�} t�EP�MQ�UR�s6����_^[���   ;���:����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HH�Qx�҃�;��:��_^[���   ;��:����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�j h�  �M��VX��_^[���   ;��:����]���������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HH�Q|�҃�;��9��_^[���   ;��9����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�j h(  �M��vW��_^[���   ;��>9����]���������������������������U����   SVWQ��4����3   ������Y�M�h(  �M���$��_^[���   ;���8����]�����������������������������U����   SVWQ��4����3   ������Y�M�j h�  �M��V��_^[���   ;��~8����]���������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E���U���Z4��_^[���   ;���7����]� �����������������������U����   SVWQ��4����3   ������Y�M��E�� %�����_^[��]��������������������������U����   SVWQ��4����3   ������Y�M��E���U���E��_^[���   ;��-7����]� �����������������������U����   SVWQ��4����3   ������Y�M��E�� %   ������_^[��]����������������������U����   SVWQ��0����4   ������Y�M��E��x ~�M��	��2����0����
ǅ0���������0���_^[���   ;��b6����]�������������������������������U����   SVWQ��4����3   ������Y�M��M��ZP���E�� hT�E�_^[���   ;���5����]����������������������U����   SVWQ��4����3   ������Y�M��E�M� +_^[��]� ��������������������������U����   SVWQ��4����3   ������Y�M��E�� tT�E�_^[��]���������������������������U����   SVWQ������=   ������Y�M��E�    �E�    �E�    �E�8 u*�MQ�M��+����uj�M���)����uǅ���    �
ǅ���   �U�������E�8 uc�M���X���} u�EP�MQ�UR�EP�MQ�M��6���7�E�E���M��rI���E��}� t�EP�MQ�UR�E�P�MQ�M���5���ыE�8 u�M��)$����tǅ���    �
ǅ���   �M�������E�8 u�M��6���EP�M���7���   �M��3X���} u�EPj �MQ�UR�EP�M��Y5���E��uh  ��=�����E�}� u3��^�M�T��P�M���@���E�E���M��H���E��}� t1�EPj �MQ�U�R�EP�M���4���Eԃ}� t�E�P�M��:O��뾋E�_^[���   ;��K3����]� �������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP��c���   �M��BH��;��|2��_^[���   ;��l2����]� ����������������������U����   SVW��@����0   �������EP�MQ�UR��c�HH���   �҃�;��
2��_^[���   ;���1����]�����������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH���   �Ѓ�;��1��_^[���   ;��1����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH���   �Ѓ�;��,1��_^[���   ;��1����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH���   �Ѓ�;��0��_^[���   ;��0����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HH���   �҃�;��E0��_^[���   ;��50����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R��c�HH���  �҃�;��/��_^[���   ;��/����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��E�� �T�E��@    �E�_^[��]�����������������U����   SVWQ��4����3   ������Y�M��M���M���E��t�E�P�"�����E�_^[���   ;���.����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� �T��E��HQ��c�Bx�H�у�;��s.��_^[���   ;��c.����]��������������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��c�Bx�H�у�;���-���} u�   �=��EP�MQ�UR�EP��c�Qx��Ѓ�;���-���M��A�E�3Ƀx ����_^[���   ;��-����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��!��E��HQ��c�Bx�H�у�;��-��_^[���   ;��-����]����������������������������U����   SVWQ������9   ������Y�M��E�P�M�Q�UR�EP�M��PP���E�;Eu�E����E�;Eu�E�����R��P��j
����XZ_^[���   ;��u,����]� �I    �j
����   �j
����   �j
l2 l1 ������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��QR��c�Hx�Q�҃�;��+��_^[���   ;��+����]� ���������������������������������������U����   SVW��@����0   �������EPQ�E�$�MQ�UR��c�HH���  �҃�;��3+��_^[���   ;��#+����]��������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��c�QH���  �Ѓ�;��*��_^[���   ;��*����]����������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP��c�QH���  �Ѓ�;��)*��_^[���   ;��*����]��������������������������������������U����   SVW��@����0   �������E,PQ�E(�$�M$Q�U R�EP�MQ�UR�EP�MQ�UR��c�HH���  �҃�(;��)��_^[���   ;��{)����]����������������������������������������U����   SVW��@����0   �������EP�MQ�UR��c�HH���  �҃�;��
)��_^[���   ;���(����]�����������������������U����   SVWQ��4����3   ������Y�M���EPQ�E�$�M�Q��c�BH���  �у�;��(��_^[���   ;��(����]� ���������������������������U����   SVWQ��(����6   ������Y�M��E�    �}u�M�����E��$�} u�M��D���E���}u�M�����E�}� u3���E�P�MQ�M���/��_^[���   ;���'����]� �����������������������������������������������U���   SVWQ�������H   ������Y�M��i"���E�}� t�} u3���   �M��)���E��}� u�E��   �E�    �	�Eԃ��EԋM�!N��9E���   �E�P�M�Q�U�R�M�$����u�̋E��E��	�Eȃ��EȋE�;E�_�Eȃ���u$�E������M������U��u��D;Du���E���P�M�����Mȃ��T��U��}��t�E�P�M�������O����E�R��P��p
����XZ_^[��   ;��k&����]� �   �p
����   �p
����   �p
b a ������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��c�Hx�Q�҃�;��%��_^[���   ;��%����]� �����������������������������������U����   SVWQ������?   ������Y�M��M��`'���E�}� u3��G  �E�    �}u�M�����E��$�} u�M���@���E���}u�M��}���E��}� u3���   �M�����E�    �	�Eԃ��EԋM����9E���   �E�P�M�����Eȃ}� u�ϋEȋHQ�M��<����t�E���P�M�����EȋHQ�M�<����t�Eԍ�   Q�M�����E����M����U�u�D;Dt&�EȋHQ�M�]<����t�Eԍ�   Q�M��I���EȋHQ�M�7<����t�Eԍ�   Q�M��#�������   _^[���   ;���#����]� ��������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B\�H0�у�;��#��_^[���   ;��#����]� �������������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP��c�QH��  �Ѓ�;��"��_^[���   ;��y"����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��  �Ѓ�;��"��_^[���   ;���!����]�������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ��c�BH���  �у�;��!��_^[���   ;��!����]������������������������������U����   SVW��@����0   ������Q�E�$Q�E�$Q���$�EP�M�D��Q�$��3�����$�MQ�M����_^[���   ;��� ����]������������������������������������U����   SVW��@����0   �������E�E������Au�E��E�E������z�E��E_^[��]���������������������������������U����   SVW������?   �����󫍍����!'��P�EP�M�Q�M�F��Q�E�$Q�E�$Q�E��$��2�����$Q�E�$Q�E�$Q�E��$�2�����$Q�E�$Q�E�$Q�E��$�2�����$�������D��P�EP�M�b9��R��P��w
���XZ_^[���   ;������]Ð   �w
����   �w
v ������������������������������������������������������������������U����   SVW��@����0   �������j �EP��c�QH��Ѓ�;�����_^[���   ;�������]��������������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;�����E�     _^[���   ;��i����]��������������������������������������U����   SVW��@����0   �������j h�  ��c�HH��҃�;����_^[���   ;�������]��������������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;�����E�     _^[���   ;��y����]��������������������������������������U����   SVW��4����3   ������h  �K'�����E��}� u3��tj �EPh�  �M���0����u�.�,j �EPh(  �M���0����u��j j�M������E��-�}� t��E�P��c�Q@�BH�Ѓ�;�����E�    3�_^[���   ;������]�������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��c���   �M��P��;����_^[���   ;������]� ����������������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;�����E�     _^[���   ;������]��������������������������������������U����   SVW��4����3   ������h�  �[%�����E��}� u3��B�EP�MQ�M�������u+�}� t��E�P��c�Q@�BH�Ѓ�;������E�    �E�_^[���   ;�������]���������������������������������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;��b���E�     _^[���   ;��I����]��������������������������������������U����   SVW��@����0   �������EP�MQ��c�BH�H�у�;�����_^[���   ;�������]�����������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;��r���E�     _^[���   ;��Y����]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH���  �у�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH���  �у�;��h��_^[���   ;��X����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH���  �Ѓ�;�����_^[���   ;�������]�������������������������U����   SVW��@����0   �������EP�MQ��c�BH���  �у�;��}��_^[���   ;��m����]��������������������������U����   SVW��@����0   �������E(P�M$Q�U R�EP�MQQ�E�$Q�E�$�UR�EP��c�QH��p  �Ѓ�$;�����_^[���   ;�������]����������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��  �Ѓ�;��l��_^[���   ;��\����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HH��  �҃�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��8  �Ѓ�;��|��_^[���   ;��l����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�QH��   �Ѓ�;�� ��_^[���   ;�������]� ��������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��$  �Ѓ�;����_^[���   ;��|����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��(  �Ѓ�;����_^[���   ;������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH��0  �у�;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH��4  �у�;��(��_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVWQ��4����3   ������Y�M�_^[��]�����������������������U����   SVW��@����0   �����󫡨c�HH��  ��;��9��_^[���   ;��)����]����������������������U����   SVW��@����0   �������EP��c�QH��  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M���E0P�M,Q�U(R�E$P�M Q�UR�EP�MQ�UR�EP�MQ�U�R��c�HH��  �҃�0;��1��_^[���   ;��!����]�, �������������������������������������������U����   SVWQ��4����3   ������Y�M���E0P�M,Q�U(R�E$P�M Q�UR�EP�MQ�UR�EP�MQ�U�R��c�HH��x  �҃�0;����_^[���   ;��q����]�, �������������������������������������������U����   SVWQ��4����3   ������Y�M���E0P�M,Q�U(R�E$P�M Q�UR�EP�MQ�UR�EP�MQ�U�R��c�HH��  �҃�0;�����_^[���   ;�������]�, �������������������������������������������U����   SVWQ��4����3   ������Y�M���E0P�M,Q�U(R�E$P�M Q�UR�EP�MQ�UR�EP�MQ�U�R��c�HH��|  �҃�0;��!��_^[���   ;������]�, �������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH��X  �Ѓ�;����_^[���   ;������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH���  �у�;��(��_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH���  �Ѓ�;����_^[���   ;������]�������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ��c�BH��\  �у�;��1��_^[���   ;��!����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR��c�HH��d  �҃�;����_^[���   ;������]���������������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U���  SVWQ��T����k   ������Y�M��}t
�   �  �M�������EP�M���M��Bp��;������E��}� u
�   �g  �EP�M�-���E���|���P�M�Z��j/��h���P�84����j��T���P�'4�����E�    �	�E����E��}��  �}� u��T���P�M�	�����h���P�M�����E�    �	�E���E�E�;E���   �E�3�;E���;M�t�ً�E�P�MQ��X���R�E���M��Bt��;������M̋P�UЋ@�E��E���T����u둍�|���P�M��]��j�E�P�M����E�P��|���QQ���$Q���$Q���$��l����/��P������R�"����P�M������.���������   R��P�،
�����XZ_^[�Ĭ  ;��P
����]� ��   ��
����   �
|���0   �
h���   �
T���   �
col2 col1 mg p �������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��4����3   ������E�@�M�	�U�B�E�@ �M�I���U�B,�E�H��ٝ<���م<���Q�$�M�A�U�
�E�@�M�A�U�J���E�@(�M�I��ٝ8���م8���Q�$�U�B�E��M��U�B�E�H���M�A$�U�J��ٝ4���م4���Q�$�M�-���E_^[���   ;������]��������������������������������������������������������������U����   SVWQ������<   ������Y�M��E�@�M��	�U��E�@�M��I���U�B$�E��H���]�E�@�M��	�U�B�E�@�M��I���U�B(�E��H���]��E�@�M��	�U�B�E�@ �M��I���U�B,�E��H���]ԋE��E���E��E��X�E��E��X�E�_^[��]� ��������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH��L  �у�;�����_^[���   ;�������]� ����������������������������������U���  SVWQ�������A   ������Y�M���E�P�� ���Q��c�Bp�Hx�у�;��h���   ���}�E_^[��  ;��I����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�Bp�H,�у�;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�Hp�QT�҃�;��X��_^[���   ;��H����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�Hp�QX�҃�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M�Q���$�M����E_^[���   ;��\����]� ����������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U���X  SVWQ�������V   ������Y�M��E��t�����   �E�P�M�))���E������M��\
���E�    �	�E����E���EP�M���M��Bp��;��F��9E���   ��E�P�MQ������R�E���M��Bt��;������M��P�U��@�E��E���T����u댋EP�MQ�U�R�E�P������Q������P�M�)����t�E��E��E��u��K����E�R��P���
����XZ_^[��X  ;������]� ��   ��
����0   ��
����   ��
p mg ���������������������������������������������������������������������������������������������������U���  SVWQ�������A   ������Y�M���E�P�� ���Q��c�BH�HH�у�;�����   ���}�E_^[��  ;������]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Qp�B(�Ѓ�;��#��_^[���   ;������]� �����������������������������U����   SVWQ������>   ������Y�M�j �M�����������EP�MQ�U�R������������Bt��;�� ���E�P�MQ�����R���������̋��P�Q�@�A�MQ�UR�E���M��Bx��;��K ���   R��P��
����XZ_^[���   ;��% ����]� �I    �
����   �
p ����������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B@�Ht�у�;��{���_^[���   ;��k�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]�  ���������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVW��@����0   ������j �EPj �MQ�UR�EP�MQ�UR�y����� _^[���   ;��������]���������������������������U����  SVW��(����v   ������ǅ���    �E�    �M�
������  �M��u����M��4�������   �EP��<�����������j h�T�������O��������P��`����t�������j j���<���Q��`���R������P�����������P������Q�1"���������P������R�"��������� P�M��h�����������uǅ(���   �
ǅ(���    ��(�����3���������� t�����ߍ������*����������t��������������������t������������������������t��������`���������������t����������������������t��������<���������3�����t.j �E,P�M�����P�MQ�UR�EP�MQ�UR�A����� �E��M���	���'j �E,Pj �MQ�UR�EP�MQ�UR������ �E��E�������M���������R��P�̜
�����XZ_^[���  ;��Z�����]Ë�   Ԝ
����   ��
����   �
_$ArrayPad icon1 �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����  SVW������z   ������M�����tj �EP�MQ��������u3��   j h   ������P�������E$P�MQ�U R�EP�MQ������R��   ���E�c��E��t�E����E�� t�E�t��E%�   t�E����E��t�E���h   ������P�MQ�URj�����R��P���
�����XZ_^[���  ;��l�����]�   ��
����   ̞
np ���������������������������������������������������������������������������������U����   SVW��@����0   ������EP�MQ�UR�EP�MQ�UR�;�����E�M���   �Eǀ�   ,��Eǀ�   ܲ�Eǀ�   ���Eǀ�   ���Eǀ�   ���Eǀ�   ��Eǀ�   w�_^[���   ;��K�����]��������������������������������������������������������U����   SVWQ��4����3   ������Y�M��8����M���E�_^[���   ;��������]�����������������������������U����   SVWQ��4����3   ������Y�M��E�P�N������E��     _^[���   ;��h�����]���������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]�����������������̋�`L����������̋�`\����������̋�`l����������̋�`@����������̋�`P����������̋�``����������̋�`D����������̋�`T����������̋�`d����������̋�`H����������̋�`X����������̋�`h�����������U����   SVWQ��4����3   ������Y�M��E�� �T�E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��M��[���E��t�E�P�������E�_^[���   ;��n�����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� �T_^[��]��������������U����   SVWQ������:   ������Y�M��E���,�����,����� ����� ��� t%��j�� ������ ������;�����������
ǅ���    _^[���   ;�������]���������������������������������������������U����   SVWQ��4����3   ������Y�M���c�P��M���l  ��;��!���_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M���c�P��M���x  ��;�����_^[���   ;�������]������������������������������U����   SVWQ������<   ������Y�M������P��c�Q�M���p  ��;��9���P�M���������������E_^[���   ;�������]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M���c�P��M���t  ��;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ��c�B��d  �у�;��-���_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP��c�Q��  �Ѓ�;������_^[���   ;�������]������������������������������U����   SVW��@����0   �����󫡨c�H��h  ��;��Y���_^[���   ;��I�����]����������������������U����   SVW��@����0   �������EP�MQ�UR��c�H��<  �҃�;������_^[���   ;��������]�����������������������U����   SVW��@����0   �������EP�MQ��c�B���  �у�;��}���_^[���   ;��m�����]��������������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVWQ������9   ������Y�M���EP�M�Q��c�B�HP�у�;������E�}� u3��x��h�T��B��P�M��Q��c�B��H  �у�;��\����E��}� u3��9��EP�M��Q�U�R�E�P��c�Q�BT�Ѓ�;��"����E�E��  �E�_^[���   ;�������]� ����������������������������������������������������������������U����   SVW������:   ������XD3ŉE��M��������EP��c�Q�BD�Ѓ�;��r����E܃}� t�E�P�M�����E�P�������E�P�M�G����M�����ER��P��
����XZ_^[�M�3�������   ;�������]ÍI     �
����   :�
����   8�
s str ������������������������������������������������������������������U����   SVW��$����7   ������XD3ŉE��M�������E�P�MQ�UR��c�H�Q|�҃�;��K����E�P�M�A����M�����ER��P��
����XZ_^[�M�3�������   ;��	�����]Ð   $�
����   0�
str ������������������������������������������������������������U����   SVW������:   ������XD3ŉE��M��������EP�MQ�UR�EPQ�E�$��c�Q�B@�Ѓ�;��N����E܃}� t�E�P�M��x���E�P�r������E�P�M�#����M�����ER��P�<�
�x���XZ_^[�M�3��e �����   ;��������]ÍI    D�
����   ^�
����   \�
s str ��������������������������������������������������������������U����   SVW��@����0   ������j h�  h�c�M������c_^[���   ;��9�����]����������������������U����   SVW��@����0   ������j h�  h�c�M�k����c_^[���   ;��������]����������������������U����   SVW��(����6   ������j h�  h�c��,���P�M�f�����������,���������c_^[���   ;��`�����]�����������������������������U����   SVW��(����6   ������j h�  h�c��,���P�M��������}����,����d����c_^[���   ;��������]�����������������������������U���  SVW�������B   ������XD3ŉE��E�E��E�    �E��D�0�Mԃ��MԋE��D�x�Mԃ��M��E�   �	�Eȃ��Eȃ}� |D�E�M������E��}�
s�E���0�MԈD��Uԃ��U���E���7�MԈD��Uԃ��U�뭋E��D� j �E�P�M������ER��P�\�
�V���XZ_^[�M�3��C�����  ;��������]Ð   d�
����   p�
hexstring ����������������������������������������������������������������������U���  SVW��t����c   ������} ��   �}   @��   j hU����������Pj0j jj �E�U�������x�����|���߭x����5Uٝt���مt���Q�$������P������P�MQ��������������!��������������E�r  �!  �} ��   �}   ��   j hU�������m���Pj0j jj �E�U�
�c�����x�����|���߭x����5Uٝt���مt���Q�$������P�������P�MQ�!������������y����������n����E��   �|�} |v	�}   vkj hU�����������Pj0j jj �m�5Uٝ|���م|���Q�$������P�\�����P�MQ�����������������������������E�Lj h U������e���P�EP��,���Q�5����P�UR�R�������,�����������������E_^[�Č  ;�������]����������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �����󫡨c�H8����;��M���_^[���   ;��=�����]��������������������������U����   SVW��@����0   �������E�Q��c�B8�H�у�;�������E�     _^[���   ;��������]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H8�Q�҃�;��X���_^[���   ;��H�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR�E�P��c�Q8�B�Ѓ�;������_^[���   ;�������]� ���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H8�Q�҃�;��H���_^[���   ;��8�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R��c�H8�Q�҃�;�����_^[���   ;�������]� ��������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��c�Q���  �Ѓ�;��5���_^[���   ;��%�����]����������������������������������U����   SVW��@����0   �������EP�MQ��c�B���  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ��c�B���  �у�;��M���_^[���   ;��=�����]��������������������������U����   SVW��@����0   �������EP�MQ��c�B���  �у�;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;��q���_^[���   ;��a�����]������������������������������U����   SVW��@����0   �������EP��c�Q�B0�Ѓ�;�����_^[���   ;��������]���������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR��c�H�Q4�҃�;�����_^[���   ;��q�����]������������������������������U����   SVW��$����7   ������XD3ŉE��M��^�����E�P��c�Q�B<�Ѓ�;������E�P�M������M��]����ER��P�d�
�M���XZ_^[�M�3��:������   ;��������]�   l�
����   x�
str ����������������������������������������������������U����   SVW��@����0   �����󫡨c�H��Q@��;��<���_^[���   ;��,�����]�������������������������U����   SVW��@����0   �������EP�MQ��c�B�HD�у�;������_^[���   ;��������]�����������������������������U����   SVW��@����0   �����󫡨c�H��QH��;��l���_^[���   ;��\�����]�������������������������U����   SVW��@����0   �����󫡨c�H��QL��;�����_^[���   ;��������]�������������������������U����   SVW��@����0   �������EP�MQ�UR��c�H�QP�҃�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP��c�Q�BT�Ѓ�;��4���_^[���   ;��$�����]���������������������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;������_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP��c�Q��|  �Ѓ�;��Q���_^[���   ;��A�����]������������������������������U����   SVW��@����0   ������E��P��P�M��@Q�U��0R�E�� P�M��Q�UR�EP��c�Q���   �Ѓ�;�����_^[���   ;�������]���������������������������������������U����   SVW��@����0   �����󫡨c�H���   ��;��I���_^[���   ;��9�����]����������������������U����   SVW��@����0   �����󫡨c�H��   ��;������_^[���   ;��������]����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQhH&  ��c�B���   �у�;��l���_^[���   ;��\�����]�����������������������������������������U����   SVW��@����0   �������EP��c�Q�B�Ѓ�;������_^[���   ;��������]���������������������������������U����   SVW������=   ������XD3ŉE��EPj h U���������P�M�Q������������������E�P��c�Q�B�Ѓ�;��L����M�����R��P��
����XZ_^[�M�3��������   ;�������]Ð   �
����    �
s ��������������������������������������������������������������U����   SVW��@����0   �������EP��c�Q�Bd�Ѓ�;�����_^[���   ;��t�����]���������������������������������U����   SVW��@����0   �������EP��c�Q�Bh�Ѓ�;�����_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP��c�Q�Bl�Ѓ�;�����_^[���   ;�������]���������������������������������U����   SVW��@����0   �����󫡨c�H��Qp��;��<���_^[���   ;��,�����]�������������������������U����   SVW��@����0   �����󫡨c�H��Qt��;������_^[���   ;��������]�������������������������U����   SVW��@����0   �����󫡨c�H��Qx��;��|���_^[���   ;��l�����]�������������������������U����   SVW��@����0   �������EP��c�Q�B|�Ѓ�;�����_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP��c�Q���   �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�UR��c�H���   �҃�;��*���_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;������_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��c�Q��X  �Ѓ�;��E���_^[���   ;��5�����]����������������������������������U����   SVW��@����0   �������EP�MQ��c�B���   �у�;������_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ��c�B���  �у�;��]���_^[���   ;��M�����]��������������������������U����   SVW������:   ������XD3ŉE��M�������E�P�MQ��c�B���   �у�;�������E�P�M�]����M��d����ER��P���
�&���XZ_^[�M�3��������   ;�������]Ð   ��
����   ��
fn ���������������������������������������������U����   SVW��@����0   �������EP�MQ��c�B���   �у�;�����_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP�MQ��c�B���  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��c�Q���  �Ѓ�;��%���_^[���   ;�������]����������������������������������U����   SVW��@����0   �������EP�MQ�UR��c�H���  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �����󫡨c�H�􋑠   ��;��I���_^[���   ;��9�����]����������������������U����   SVW��@����0   �������EP�MQ��c�B���  �у�;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP��c�Q��P  �Ѓ�;��q���_^[���   ;��a�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR��c�H��T  �҃�;������_^[���   ;��������]�����������������������U����   SVW�� ����8   ������XD3ŉE��M��c�����E�P��c�Q���   �Ѓ�;������E�P�M�����M�������ER��P���
�ʿ��XZ_^[�M�3��������   ;��=�����]Ð   ��
����   ��
bc �������������������������������������������������U����   SVW��@����0   �����󫡨c�H�􋑰  ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   �������EP��c�Q��\  �Ѓ�;��Q���_^[���   ;��A�����]������������������������������U����   SVW��,����5   �������EP��0���Q��c�B���   �у�;�������U��
�H�J�@�B�E_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP�MQ��c�B��  �у�;��M���_^[���   ;��=�����]��������������������������U����   SVW��@����0   �������EPQ�E�$Q�E�$�MQ��c�B���   �у�;������_^[���   ;�������]����������������������������U����   SVW��@����0   �������EP�MQ�UR��c�H���   �҃�;��Z���_^[���   ;��J�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR��c�H��   �҃�;������_^[���   ;��������]�����������������������U����   SVW��@����0   �������EP�MQ�UR��c�H��  �҃�;��z���_^[���   ;��j�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR��c�H���  �҃�;��
���_^[���   ;��������]�����������������������U����   SVW��@����0   �������EP�MQ�UR��c�H��$  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ��c�B��(  �у�;��-���_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ��c�B��,  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP��c�Q��0  �Ѓ�;��Q���_^[���   ;��A�����]������������������������������U����   SVW��@����0   �������EP��c�Q��4  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP��c�Q��8  �Ѓ�;��q���_^[���   ;��a�����]������������������������������U����   SVW��@����0   �������EP��c�Q��<  �Ѓ�;�����_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP��c�Q��@  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P��c�Q��D  �Ѓ�;�������u3���E�R��P�@�
�g���XZ_^[���   ;��������]�   H�
����   x�
����   q�
����   l�
data sub_id main_id ������������������������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P��c�Q��D  �Ѓ�;�� �����u3���E�R��P�0�
�w���XZ_^[���   ;��������]�   8�
����   h�
����   a�
����   \�
data sub_id main_id ������������������������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P��c�Q��D  �Ѓ�;��0�����u3���E�R��P� �
臵��XZ_^[���   ;�������]�   (�
����   X�
����   Q�
����   L�
data sub_id main_id ������������������������������������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;��Q���_^[���   ;��A�����]������������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M�����P�U�R��c�H0���   �҃�(;�����_^[���   ;�������]�$ ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M����P�U�R��c�H0���   �҃�(;��Ŀ��_^[���   ;�贿����]�$ ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P��c�Q0���   �Ѓ�(;��ؾ��_^[���   ;��Ⱦ����]�$ ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��c�B0���   �у�;��L���_^[���   ;��<�����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q0���   �Ѓ�;��̽��_^[���   ;�輽����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H0���   �҃�;��U���_^[���   ;��E�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��c�B0���   �у�;��̼��_^[���   ;�輼����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q0���   �Ѓ�;��L���_^[���   ;��<�����]�������������������������U����   SVW��@����0   �����󫡨c�H0�􋑼   ��;�����_^[���   ;��ٻ����]����������������������U����   SVW��@����0   �������E�Q��c�B0���   �у�;������E�     _^[���   ;��f�����]�����������������������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;�葺��_^[���   ;�聺����]������������������������������U����   SVW��@����0   �����󫡨c�H���  ��;��)���_^[���   ;�������]����������������������U����   SVW��@����0   �����󫡨c�H��  ��;��ɹ��_^[���   ;�蹹����]����������������������U����   SVW��@����0   �������EP��c�Q��,  �Ѓ�;��a���_^[���   ;��Q�����]������������������������������U����   SVW��@����0   �������EP��c�Q��8  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP��c�Q��0  �Ѓ�;�聸��_^[���   ;��q�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��c�Q��(  �Ѓ�;�����_^[���   ;��������]����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ��c�B��H  �у�;�職��_^[���   ;��q�����]������������������������������U����   SVW��0����4   �������EP�MQ�UR��4���P��c�Q���  �Ѓ�;�����P�M�l�����4����J����E_^[���   ;��۶����]����������������������������������������U����   SVW������;   ������j hLGOg���������PhicMC�E�P������������蹦���M��ʫ����u�M�����M������E��M�詫��P�M������M������ER��P� �
舩��XZ_^[���   ;�������]Ð   (�
����   4�
dat ��������������������������������������������������������U����   SVW��@����0   �������EP�MQ��c�B��`  �у�;��m���_^[���   ;��]�����]��������������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW������9   ������EP��MQ�� ���R��c�H���  �҃�;�致�����_����� ��������E_^[���   ;��b�����]�������������������������������U����   SVW��@����0   �������EP�MQ��c�B���  �у�;������_^[���   ;�������]��������������������������U����   SVW��(����6   �������EP��,���Q��c�B���  �у�;�芳��P�M������,���������E_^[���   ;��c�����]��������������������������������U����   SVW��(����6   �������EP��,���Q��c�B���  �у�;������P�M������,����U����E_^[���   ;��Ӳ����]��������������������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;��q���_^[���   ;��a�����]������������������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP��c�Q��   �Ѓ�;�葱��_^[���   ;�聱����]������������������������������U����   SVW��@����0   �������E$P�M Q�UR�EP�MQ�UR�EP�MQ��c�B��  �у� ;�����_^[���   ;��������]����������������������������������U����   SVW��@����0   �������E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR��c�H��  �҃�$;��r���_^[���   ;��b�����]�������������������������������U����   SVW������9   ������EP�MQ�UR���̋EP�{�����,���Q��c�B���  �у�P�M������,����H����E_^[���   ;��Ư����]�����������������������������������U����   SVW��0����4   �������EP�MQ�UR��4���P��c�Q��  �Ѓ�;��R���P�M輯����4���蚼���E_^[���   ;��+�����]����������������������������������������U����  SVW��(����6  ������XD3ŉE��E�E�E�P�MQ������R�B�����������Ph$U��c�Q���  �Ѓ�;�蒮���E�    R��P���
����XZ_^[�M�3���������  ;��`�����]�   ��
����   ��
t ������������������������������������������������������U����   SVW��(����6   �������,���P��c�Q��h  �Ѓ�;��έ��P�M�Ǻ����,����)����E_^[���   ;�觭����]������������������������������������U����   SVW��(����6   �������,���P��c�Q��l  �Ѓ�;��>���P�M�7�����,��������E_^[���   ;�������]������������������������������������U����   SVW������<   ������XD3ŉE��S�����u�\h���M������EPh���M������EPh���M�����j �E�PhicMC�����Q������������Ź���M�跜��R��P���
�ß��XZ_^[�M�3��������   ;��6�����]Ë�   ��
����   �
msg ��������������������������������������������������������U����   SVW������<   ������XD3ŉE��C�����u�M�����E�^h!���M������EPh!���M�����j �E�PhicMC�����Q����������T���P�M�\��������諸���M�蝛���ER��P��
覞��XZ_^[�M�3��������   ;�������]Ð   �
����    �
msg ������������������������������������������������������������U����   SVW������?   ������XD3ŉE��#�����u3��^h#���M������EPh#���M��h���j �E�PhicMC�����Q���������>�������������藷���M�艚�������R��P�$�
菝��XZ_^[�M�3��|������   ;�������]Ë�   ,�
����   8�
msg ��������������������������������������������������������������������U����   SVW������?   ������XD3ŉE�������u3��^hs���M��l����EPhs���M��H���j �E�PhicMC�����Q������������������������w����M��i��������R��P�D�
�o���XZ_^[�M�3��\������   ;�������]Ë�   L�
����   X�
msg ��������������������������������������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR��c�H��,  �҃�;��.���_^[���   ;�������]���������������������������U����   SVW��@����0   �������EP�MQ�UR��c�H���  �҃�;�躧��_^[���   ;�誧����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR��c�H��0  �҃�;��>���_^[���   ;��.�����]���������������������������U����   SVW��@����0   ������E�8 t#��E�Q��c�B���  �у�;��Ǧ���E�     _^[���   ;�讦����]���������������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;��Q���_^[���   ;��A�����]������������������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;�����_^[���   ;��ѥ����]������������������������������U����   SVW��@����0   �������EP�MQ�UR��c�H���  �҃�;��j���_^[���   ;��Z�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR��c�H���  �҃�;������_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR��c�H���  �҃�;�芤��_^[���   ;��z�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR��c�H���  �҃�;�����_^[���   ;��
�����]�����������������������U����   SVW��@����0   �����󫡨c�H���  ��;�蹣��_^[���   ;�詣����]����������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP��c�Q���  �Ѓ�;��9���_^[���   ;��)�����]��������������������������������������U����   SVW��@����0   �������EP�MQ��c�B���  �у�;�轢��_^[���   ;�譢����]��������������������������U����   SVW��@����0   �����󫡨c�H���  ��;��Y���_^[���   ;��I�����]����������������������U����   SVW��$����7   �������EP��(���Q��c�B���  �у�;�����P�M�q�����(����,����E_^[���   ;��á����]��������������������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;��a���_^[���   ;��Q�����]������������������������������U����   SVW��@����0   �������EP��c�Q��   �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ��c�B��  �у�;��}���_^[���   ;��m�����]��������������������������U����   SVW��@����0   �������EP��c�Q��  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�UR��c�H��  �҃�;�蚟��_^[���   ;�芟����]�����������������������U����   SVW��@����0   �������EP�MQ�UR��c�H��  �҃�;��*���_^[���   ;�������]�����������������������U����   SVW������;   ������h������������j �����PhicMC��4���Q�C�������4�����������������_^[���   ;�菞����]��������������������������������������������U����   SVW��@����0   �������EP�MQ�UR��c�H��   �҃�;�����_^[���   ;��
�����]�����������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;�豝��_^[���   ;�衝����]������������������������������U����   SVW��@����0   �������EP�MQ�UR��c�H��L  �҃�;��:���_^[���   ;��*�����]�����������������������U����   SVW��@����0   �����󫡨c�H��P  ��;��ٜ��_^[���   ;��ɜ����]����������������������U����   SVW��@����0   �������EP�MQ�UR��c�H��T  �҃�;��j���_^[���   ;��Z�����]�����������������������U����   SVW��4����3   ������j �M�݋���E��}� t�E�P襝�����E�P�i�����R��P�P�
�Y���XZ_^[���   ;��֛����]Ë�   X�
����   d�
c ������������������������������������������U����   SVW��@����0   �����󫡨c�H$��Q��;��\���_^[���   ;��L�����]�������������������������U����   SVW��@����0   �������EP��c�Q$�B�Ѓ�;������_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP��c�Q$�B�Ѓ�;�脚��_^[���   ;��t�����]���������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q$�BD�Ѓ�;������E�_^[���   ;��������]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q$�BD�Ѓ�;�蟙����EP�M�Q��c�B$�Hd�у�;��}����E�_^[���   ;��j�����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q$�BD�Ѓ�;��������EP�M�Q��c�B$�H�у�;��ݘ���E�_^[���   ;��ʘ����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q$�BD�Ѓ�;��_�����E�P�MQ��c�B$�HL�у�;��=����E�_^[���   ;��*�����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q$�BH�Ѓ�;�迗��_^[���   ;�诗����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B$�HL�у�;��K���_^[���   ;��;�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q$�B�Ѓ�;��ϖ��_^[���   ;�迖����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q$�B�Ѓ�;��S���_^[���   ;��C�����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q$�B�Ѓ�;��ӕ��_^[���   ;��Õ����]� �����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q$�B�Ѓ�;��_���_^[���   ;��O�����]����������������������������U����   SVWQ������=   ������Y�XD3ŉE��M�M��9�����E�P��c�Q$�B�Ѓ�;��ݔ���EЃ}� t�E�P�M��\����E�P�������E�P�M財���M������ER��P������XZ_^[�M�3���������   ;��z�����]�    �����   �����   �str s ��������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�Hp�у�;��˓��_^[���   ;�軓����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B$�H�у�;��K���_^[���   ;��;�����]� �������������������������������������U���   SVWQ�� ����@   ������Y�XD3ŉE��M�M��l�����E�P��c�Q$�B �Ѓ�;�轒���Eă}� t�E�P�M��J����E�P�������E�P�M�����M��%����ER��P������XZ_^[�M�3��ԧ����   ;��Z�����]�    �����   �����   �fn f ���������������������������������������������������������������U���   SVWQ�� ����@   ������Y�XD3ŉE��M�M��L�����E�P��c�Q$�B$�Ѓ�;�蝑���Eă}� t�E�P�M��*����E�P��������E�P�M������M������ER��P���Ǆ��XZ_^[�M�3�账����   ;��:�����]�    �����   ����   fn f ���������������������������������������������������������������U����   SVWQ������<   ������Y�M��EP�����Q�M��m������r��������%����E_^[���   ;��u�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q$�B(�Ѓ�;�����_^[���   ;��������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q$�Bh�Ѓ�;�蟏��_^[���   ;�菏����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B$�H,�у�;��+���_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B$�H0�у�;�諎��_^[���   ;�蛎����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B$�H4�у�;��+���_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B$�H8�у�;�諍��_^[���   ;�蛍����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ��c�B$�HL�у�;��+����E�_^[���   ;�������]� ����������������������������������U����   SVW������:   ������XD3ŉE��EP�M��J�����EP�M�Q��c�B$�H@�у�;�蚌���E�P�M�����M��#����ER��P��
����XZ_^[�M�3��ҡ�����   ;��X�����]�   �
����   �
fn ���������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B$�H@�у�;��ˋ���E�_^[���   ;�踋����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B$�H<�у�;��K���_^[���   ;��;�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B$�H<�у�;��ˊ�������_^[���   ;�贊����]� ������������������������������U����   SVW��@����0   ������E�8 t ��E�Q��c�B$�H�у�;��J����E�     _^[���   ;��1�����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H$�QP�҃�;��ȉ��_^[���   ;�踉����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B$�HT�у�;��K���_^[���   ;��;�����]� �������������������������������������U����   SVW��@����0   �����󫡨c�H$��QX��;��܈��_^[���   ;��̈����]�������������������������U����   SVW��@����0   �������EP��c�Q$�B\�Ѓ�;��t���_^[���   ;��d�����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q$�B`�Ѓ�;�����_^[���   ;�������]� �����������������������������U����   SVW��@����0   �����󫡨c�H(����;�荇��_^[���   ;��}�����]��������������������������U����   SVW��@����0   �������E�Q��c�B(�H�у�;��"����E�     _^[���   ;��	�����]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR�E�P��c�Q(�B�Ѓ�;�臆��_^[���   ;��w�����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q(�B�Ѓ�;�����_^[���   ;��������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B(�H�у�;�蛅��_^[���   ;�苅����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q(�B�Ѓ�;�����_^[���   ;�������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H(�Q�҃�;�蘄��_^[���   ;�舄����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���j�EP�MQ�U�R��c�H(�Q�҃�;�����_^[���   ;�������]� ��������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H(�Q�҃�;�蘃��_^[���   ;�舃����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q(�B �Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q(�B$�Ѓ�;�诂��_^[���   ;�蟂����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q(�B(�Ѓ�;��?���_^[���   ;��/�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B(�H,�у�;��ˁ��_^[���   ;�軁����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B(�HP�у�;��K���_^[���   ;��;�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B(�HT�у�;��ˀ��_^[���   ;�軀����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B(�HX�у�;��K���_^[���   ;��;�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B(�H\�у�;�����_^[���   ;������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B(�H`�у�;��K��_^[���   ;��;����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B(�Hp�у�;���~��_^[���   ;��~����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B(�Hd�у�;��K~��_^[���   ;��;~����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B(�Hh�у�;���}��_^[���   ;��}����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B(�Hl�у�;��K}��_^[���   ;��;}����]� �������������������������������������U����   SVWQ������?   ������Y�M��E�    �E�    �E�P�M��i����u3���   �}� u)����������P�M��������������   �   ��h(U��B��P�M�Q��c�B��H  �у�;��j|���E��}� uj��M��B���3��Lj �E�P�M�Q�M�舔����u�E�P�v����3��&j �E��P�M�Q�M譠���E�P�~v�����   R��P�@�io��XZ_^[���   ;���{����]�    H����   b����   `c len ������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q�Bd�Ѓ�;��{��_^[���   ;��{����]� �����������������������������U���   SVWQ�� ����@   ������Y�XD3ŉE��M�M������E�P�M��u����uǅ���    �M������������$�E�P�M�i��ǅ���   �M��Ғ�������R��P���m��XZ_^[�M�3�謏����   ;��2z����]�    �����   str ����������������������������������������������������U����   SVWQ��(����6   ������Y�M��E�P�M��p����u3���E�����؋M��   R��P����l��XZ_^[���   ;��ty����]� ��   �����   �c ��������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��+�����t�M��Q�M�������tǅ0���   �
ǅ0���    ��0���_^[���   ;��x����]� ����������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M�苏����t2�M��Q�M��x�����t�U��R�M��e�����tǅ0���   �
ǅ0���    ��0���_^[���   ;��x����]� �������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��^�����t2�M��Q�M��K�����t�U��R�M��8�����tǅ0���   �
ǅ0���    ��0���_^[���   ;��[w����]� �������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��]a����tE�M��Q�M��Ja����t2�U��R�M��7a����t�E��$P�M��$a����tǅ0���   �
ǅ0���    ��0���_^[���   ;��v����]� ��������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��a����tE�M��Q�M��ya����t2�U��0R�M��fa����t�E��HP�M��Sa����tǅ0���   �
ǅ0���    ��0���_^[���   ;���u����]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M��} ����Q�M�茄��_^[���   ;��Ju����]� ��������������������U����   SVWQ��0����4   ������Y�M��EQ� �$�M��Tm����t"�MQ�A�$�M��>m����tǅ0���   �
ǅ0���    ��0���_^[���   ;��t����]� ��������������������������������U����   SVWQ��0����4   ������Y�M��EQ� �$�M��l����t8�MQ�A�$�M��l����t"�UQ�B�$�M��l����tǅ0���   �
ǅ0���    ��0���_^[���   ;�� t����]� ������������������������������������������U����   SVWQ��0����4   ������Y�M��E��� �$�M��Ji����t<�M���A�$�M��2i����t$�U���B�$�M��i����tǅ0���   �
ǅ0���    ��0���_^[���   ;��:s����]� ����������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��\����tE�M��Q�M���[����t2�U��R�M���[����t�E��$P�M���[����tǅ0���   �
ǅ0���    ��0���_^[���   ;��hr����]� ��������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M�������tE�M��Q�M�������t2�U��0R�M�������t�E��HP�M��ہ����tǅ0���   �
ǅ0���    ��0���_^[���   ;��q����]� ��������������������������������������������������U����   SVWQ������=   ������Y�M�j �M�h�����E���h(U��B��P�M�Q��c�B��H  �у�;���p���Eԃ}� uj��M��֔��3��dj �E�P�M�Q�M�R����E�P�M��܊����t �M�Q�U�R�M���{����tǅ���   �
ǅ���    ������E�E�P��j�����E�R��P��&��c��XZ_^[���   ;��bp����]�    �&����   �&mem ������������������������������������������������������������������������������������U����   SVWQ������<   ������Y�M��� ���P�M�^��P�M�蚀��������� ������������_^[���   ;��o����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M����EP�M�Q��c�B(�H0�у�;��o��_^[���   ;��
o����]� ������������������������������������U����   SVWQ��4����3   ������Y�M����EP�M�Q��c�B(�H4�у�;��n��_^[���   ;��n����]� ������������������������������������U����   SVWQ��4����3   ������Y�M����EP�M�Q��c�B(�H8�у�;��n��_^[���   ;��
n����]� ������������������������������������U����   SVWQ��4����3   ������Y�M����EP�M�Q��c�B(�H<�у�;��m��_^[���   ;��m����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B(�H@�у�;��m��_^[���   ;��m����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H(�Qt�҃�;��l��_^[���   ;��l����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B(�HD�у�;��l��_^[���   ;��l����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$�E�P��c�Q(�BH�Ѓ�;��k��_^[���   ;��k����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�E�P��c�Q(�BL�Ѓ�;��k��_^[���   ;��k����]� ��������������������������������U����   SVW��@����0   �����󫡨c�H,��Q��;��j��_^[���   ;��j����]�������������������������U����   SVWQ��4����3   ������Y�M���c�P,��M��B8��;��Dj��_^[���   ;��4j����]���������������������������������U����   SVW��@����0   �������E�Q��c�B,�H �у�;���i���E�     _^[���   ;��i����]��������������������������������������U����   SVWQ��4����3   ������Y�M���c�P,��M��B<��;��Ti��_^[���   ;��Di����]���������������������������������U����   SVWQ������<   ������Y�M������P��c�Q,�M��B@��;���h��P�M�av��������e]���E_^[���   ;��h����]� �������������������������������U����   SVWQ������9   ������Y�M���EP�� ���Q��c�B,�M��PH��;��Hh��P�M�Au���� ���裀���E_^[���   ;��!h����]� �������������������������������������������U����   SVW��@����0   �������j j ��c�H,��҃�;��g��_^[���   ;��g����]�����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H,�Q�҃�;��8g��_^[���   ;��(g����]� ����������������������������������U����   SVW��@����0   �������E�Q��c�B,�H�у�;���f���E�     _^[���   ;��f����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q,�B�Ѓ�;��?f��_^[���   ;��/f����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q,�B�Ѓ�;���e��_^[���   ;��e����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q,�B�Ѓ�;��_e��_^[���   ;��Oe����]����������������������������U����   SVWQ��4����3   ������Y�M���c�P,��M��B,��;���d��_^[���   ;���d����]���������������������������������U����   SVWQ��4����3   ������Y�M���c�P,��M��BD��;��d��_^[���   ;��td����]���������������������������������U����   SVWQ��4����3   ������Y�M���c�P,��M��B0��;��d��_^[���   ;��d����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��c�B,�M��P4��;��c��_^[���   ;��c����]� �������������������������������������U����   SVW��@����0   �������EP�MQ�UR��c�H,�Q$�҃�;��c��_^[���   ;��c����]��������������������������U����   SVW��@����0   �������EP�MQ�UR��c�H,�QL�҃�;��b��_^[���   ;��b����]��������������������������U����   SVW��@����0   �������EP��c�Q,�B(�Ѓ�;��Db��_^[���   ;��4b����]���������������������������������U���   SVWQ�� ����@   ������Y�XD3ŉE��M�M��ll����E�P��c�Q,�B�Ѓ�;��a���Eă}� t�E�P�M��Jo���E�P�������E�P�M�o���M��%V���ER��P��5��T��XZ_^[�M�3���v����   ;��Za����]�    �5����   �5����   �5fn f ���������������������������������������������������������������U����   SVW��@����0   �������EP�MQ��c�B�H�у�;��`��_^[���   ;��`����]�����������������������������U����   SVW��@����0   �������EP�MQ�UR��c�H�Q�҃�;��=`��_^[���   ;��-`����]��������������������������U����   SVW��@����0   �������EP�MQ��c�B�H�у�;���_��_^[���   ;���_����]�����������������������������U����   SVW��@����0   �������EP�MQ�UR��c�H�Q�҃�;��]_��_^[���   ;��M_����]��������������������������U����   SVW��@����0   �������EP�MQ��c�B�H�у�;���^��_^[���   ;���^����]�����������������������������U����   SVW��@����0   �������EP�MQ��c�B��\  �у�;��}^��_^[���   ;��m^����]��������������������������U����   SVW��@����0   �������EP��c�Q�B �Ѓ�;��^��_^[���   ;��^����]���������������������������������U����   SVW��@����0   �������EP��c�Q�B$�Ѓ�;��]��_^[���   ;��]����]���������������������������������U����   SVW��@����0   �������EP�MQ��c�B�H,�у�;��0]��_^[���   ;�� ]����]�����������������������������U����   SVW������=   ������XD3ŉE��M��ag����c�H��Q(��;��\���EЃ}� t�E�P�M��Gj���E�P�|�����E�P�M�j���M��"Q���ER��P��:��O��XZ_^[�M�3���q�����   ;��W\����]ÍI    �:����   �:����   �:fn f �����������������������������������������������������������U����   SVW������=   ������XD3ŉE��M��Qf����c�H��X  ��;��[���EЃ}� t�E�P�M��4i���E�P� {�����E�P�M�i���M��P���ER��P��;��N��XZ_^[�M�3��p�����   ;��D[����]�   �;����   <����    <fn f �����������������������������������������������������������U����   SVW��@����0   �������EP�MQ��c�B��d  �у�;��Z��_^[���   ;��Z����]��������������������������U���$  SVW�������I   ������ǅ8���    �=|h t!������P�|h��M����8����������������d����8���������������������������R�M�yg����8�����t��8����������kN����8�����t��8�����������NN���E_^[��$  ;��Y����]�����������������������������������������������������������U����   SVW������9   �������EP�� ���Q��c�B��L  �у�;��Y��P�M�f���� ����M���E_^[���   ;���X����]��������������������������������U����   SVW��@����0   ������j�EP��p�����E_^[���   ;��X����]������������������������������U����   SVW��@����0   �����󫡨c�H���   ��;��9X��_^[���   ;��)X����]����������������������U����   SVW��@����0   �������EP��c�Q���   �Ѓ�;���W���E�     _^[���   ;��W����]�������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q���   �Ѓ�;��@W��_^[���   ;��0W����]� ��������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q���   �Ѓ�;���V��_^[���   ;��V����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q���   �Ѓ�;��\V��_^[���   ;��LV����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�HL�у�;���U��_^[���   ;���U����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�HP�у�;��kU��_^[���   ;��[U����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�HT�у�;���T��_^[���   ;���T����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�HX�у�;��kT��_^[���   ;��[T����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H\�у�;���S��_^[���   ;���S����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H`�у�;��kS��_^[���   ;��[S����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B���   �у�;���R��_^[���   ;���R����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�Hd�у�;��kR��_^[���   ;��[R����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�Hh�у�;���Q��_^[���   ;���Q����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�Hl�у�;��kQ��_^[���   ;��[Q����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�Hp�у�;���P��_^[���   ;���P����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�Ht�у�;��kP��_^[���   ;��[P����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�Hx�у�;���O��_^[���   ;���O����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H|�у�;��kO��_^[���   ;��[O����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B���   �у�;���N��_^[���   ;���N����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B���   �у�;��hN��_^[���   ;��XN����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B���   �у�;���M��_^[���   ;���M����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B���   �у�;��hM��_^[���   ;��XM����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H���   �҃�;���L��_^[���   ;���L����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H���   �҃�;��eL��_^[���   ;��UL����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B���   �у�;���K��_^[���   ;���K����]� ����������������������������������U����   SVWQ��0����4   ������Y�M��} t2��EP�M�Q��c�B �H(�у�;��eK����tǅ0���   �
ǅ0���    ��0���_^[���   ;��5K����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�UR��c�H �Qh�҃�;��J��_^[���   ;��J����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��} u3��'��EP�M�Q��c�B �H,�у�;��1J���   _^[���   ;��J����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M����EP�M�Q��c�B��у�;��I��_^[���   ;��I����]� �������������������������������������U����   SVWQ��4����3   ������Y�M����EP�M�Q��c�B�H�у�;��*I��_^[���   ;��I����]� ������������������������������������U����   SVWQ��4����3   ������Y�M����EP�M�Q��c�B�H�у�;��H��_^[���   ;��H����]� ������������������������������������U����   SVWQ��4����3   ������Y�M����EP�M�Q��c�B�H�у�;��*H��_^[���   ;��H����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H�у�;��G��_^[���   ;��G����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H�у�;��+G��_^[���   ;��G����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H���   �҃�;��F��_^[���   ;��F����]� �������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$�E�P��c�Q�B�Ѓ�;��(F��_^[���   ;��F����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�E�P��c�Q�B�Ѓ�;��E��_^[���   ;��E����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H �у�;��+E��_^[���   ;��E����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H$�у�;��D��_^[���   ;��D����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H(�у�;��+D��_^[���   ;��D����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H,�у�;��C��_^[���   ;��C����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H0�у�;��+C��_^[���   ;��C����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H4�у�;��B��_^[���   ;��B����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H8�у�;��+B��_^[���   ;��B����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H<�у�;��A��_^[���   ;��A����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��c�B���   �у�;��A��_^[���   ;��A����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�HD�у�;��@��_^[���   ;��@����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B���   �у�;��@��_^[���   ;��@����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H�QH�҃�;��?��_^[���   ;��?����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q���   �Ѓ�;��?��_^[���   ;��?����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B���   �у�;��>��_^[���   ;��>����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B���   �у�;��(>��_^[���   ;��>����]� ����������������������������������U����   SVWQ��4����3   ������Y�M����EP�M�Q��c�B���   �у�;��=��_^[���   ;��=����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H���   �҃�;��%=��_^[���   ;��=����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q���   �Ѓ�;��<��_^[���   ;��<����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H���   �҃�;��5<��_^[���   ;��%<����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q���   �Ѓ�;��;��_^[���   ;��;����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q���   �Ѓ�;��L;��_^[���   ;��<;����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q���   �Ѓ�;���:��_^[���   ;���:����]�������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ��c�B���   �у�;��a:��_^[���   ;��Q:����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��c�Q���   �Ѓ�;���9��_^[���   ;���9����]����������������������������������U����   SVW��(����6   �������EP�MQ��,���R��c�H��4  �҃�;��g9��P�M�`F����,�����Q���E_^[���   ;��@9����]���������������������������������������������U����   SVW��@����0   �������EP�MQ��c�B��8  �у�;���8��_^[���   ;��8����]��������������������������U���(  SVW�������J   ������XD3ŉE��E�    �M��,%���} tg��EP��c�Q4�B�Ѓ�;��E8���Ẽ}� uǅ����    �M��(����������   ��E�P�MQ�Ű�M̋P(��;��8���E��b��EP��c�Q0�B�Ѓ�;���7���E��}� uǅ����    �M��(���������j��E�P�MQ�U���M��P ��;��7���E�M��7V�����t%��E�P�MQ��c�B0���   �у�;��h7���E������M��'��������R��P� `�*��XZ_^[�M�3��L����(  ;��&7����]Ë�   `����   `result ���������������������������������������������������������������������������������������������������������������������U����   SVWQ������:   ������Y�M��M�
U������������NIVbb�����NIVb�  �����TCAb5�����TCAb��  �����$'  ��  �����MicM�.  ��  �����INIbt]�  �����atni-�����atnit6�����ckhc�Z  �����ytsdt\�  �����cnys��   �o  �+���e  �E��x t
�   �T  �E��@   �E����M��B��;��f5���/  �E����M��B��;��K5���E��@    �  �E��x u
�   ��   �E����M��B��;��5����   j hIicM�M��]���E��EP�M�Q�U���M��P��;���4���   j hIicM�M�]���E��EP�M�Q�U���M��P��;��4���uj hdiem�M�]���E��EP�M�Q�U���M��P��;��w4���E��E��=�E����M��B��;��Y4���%�!��EP�M���M��B��;��;4���   �3�_^[���   ;��"4����]� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E�� xU��E�Phߠ��c�Q0��Ѓ�;��"3���M��A�E��@    �E�_^[���   ;���2����]��������������������������������������������U����   SVWQ��4����3   ������Y�M��M��1���E��t�E�P�-&�����E�_^[���   ;��~2����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� xU�E��x t!��E��HQ��c�B0�H�у�;��
2���E��@    _^[���   ;���1����]���������������������������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��c�B0���   �у�;��y1��_^[���   ;��i1����]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��c�H0���   �҃�;���0��_^[���   ;���0����]� ��������������������������������U����   SVWQ��4����3   ������Y�M��M��-����P��c�H0���   �҃�;��x0��_^[���   ;��h0����]�������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j4�E��HQ��c�B0���   �у�(;���/��_^[���   ;���/����]������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j;�E��HQ��c�B0���   �у�(;��W/��_^[���   ;��G/����]������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��,��P��c�Q0���   �Ѓ�;���.��_^[���   ;���.����]� �����������������������������U���  SVWQ�������A   ������Y�XD3ŉE��M�E P�M���W���EPh8kds�M��QV���E�    ��E�P�M�Qj �UR�EP�MQ�UR�EPj2�M��K+��P��c�Q0���   �Ѓ�(;��	.���Ẻ� ����M��N���� ���R��P�`i�T!��XZ_^[�M�3��AC����  ;���-����]� �   hi����   �i����   �ir customdata �������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��K*����P��c�H0���   �҃�;��-��_^[���   ;���,����]�������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��t��j j j j j �E Pj �MQj�U��BP��c�Q0���   �Ѓ�(;��f,����EP�MQ�UR�EPj �MQ�U��BP��c�Q0���   �Ѓ�;��,,��_^[���   ;��,����]� ������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��!��E��HQ��c�B0�H�у�;��+��_^[���   ;��+����]����������������������������U����   SVWQ��4����3   ������Y�M��M���.��_^[���   ;��%+����]� �������������������������������U����   SVWQ��$����7   ������Y�M��E��x uj �M�Q���E�X�M�)����P�EP�M�zO��P�M��QR��(���P��c�Q0���   �Ѓ�;��*��P�M��*����(�����7���E_^[���   ;��]*����]� �������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��c�H0�Q �҃�;��Y)��_^[���   ;��I)����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��E��x u�7��j j j j j j �EPj j�M��QR��c�H0���   �҃�(;��(��_^[���   ;��(����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��6�M�'����P�EP�M�M��P�M��QR��c�H0�Q�҃�;��(��_^[���   ;��
(����]� ������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��6�M�|&����P�EP�M�eL��P�M��QR��c�H0�Ql�҃�;��z'��_^[���   ;��j'����]� ������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��_�E��ًU�
�E��ًU�
��EP�MQ�U��BP��c�Q4�Bl�Ѓ�;���&���E�E��ًU�
�E��ًU�
�E�_^[���   ;��&����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��)��EP�MQ�U��BP��c�Q4�Bl�Ѓ�;��&��_^[���   ;��&����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��)��EP�MQ�U��BP��c�Q4�Bt�Ѓ�;��%��_^[���   ;��w%����]� ���������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��_�E��ًU�
�E��ًU�
��EP�MQ�U��BP��c�Q4�Bt�Ѓ�;���$���E�E��ًU�
�E��ًU�
�E�_^[���   ;��$����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M�h���h  ��EPj 3Ƀ} ����Qj �UR�EP�M��-��_^[���   ;��$����]� ����������������������������������������U���  SVWQ�������B   ������Y�XD3ŉE��M�htniv�M���B���EPhulav�M��K��hgnlfhtmrf�M��K���EPhinim�M��}K���EPhixam�M��lK���EPhpets�M��[K���EPhsirt�M��JK���}   �u	�}$���t"�E Ph2nim�M��'K���E$Ph2xam�M��K���E�P�MQ�����R�M��W������5��������������H0���M��:��������R��P�tt�@��XZ_^[�M�3��-8����  ;��"����]�  �   |t����   �tmsg ����������������������������������������������������������������������������������������������������U���  SVWQ�������B   ������Y�XD3ŉE��M�htlfv�M��A��Q�E�$hulav�M������EPhtmrf�M���I��Q�E�$hinim�M����Q�E�$hixam�M����Q�E�$hpets�M��z���E,Phsirt�M��I���E ��.����Dz�E$��.����D{(Q�E �$h2nim�M��5��Q�E$�$h2xam�M��!���E(Phdauq�M��&I���E�P�MQ�����R�M��g������3��������������X.���M��J��������R��P�dv�P��XZ_^[�M�3��=6����  ;��� ����]�( �   lv����   xvmsg ����������������������������������������������������������������������������������������������������U����   SVWQ��0����4   ������Y�M��E$Pj Q���$Q���$haerfQ�E �$Q�E�$Q�E�$�MQ��$�UR�M�� J������   �E$Pj Q���$Q���$haerfQ�E �$Q�E�$Q�E�$�MQ�A�$�UR�M���I����tR�E$Pj Q���$Q���$haerfQ�E �$Q�E�$Q�E�$�MQ�A�$�UR�M��I����tǅ0���   �
ǅ0���    ��0���_^[���   ;������]�  ��������������������������������������������������������������������������������������U����   SVWQ��0����4   ������Y�M��E$PQ�E �$Q�E�$Q�E�$�MQ��$�UR�M��@����tr�E$PQ�E �$Q�E�$Q�E�$�MQ�A�$�UR�M���?����t?�E$PQ�E �$Q�E�$Q�E�$�MQ�A�$�UR�M��?����tǅ0���   �
ǅ0���    ��0���_^[���   ;�������]�  �������������������������������������������������������������������U����   SVWQ��0����4   ������Y�M��E$PQ�E �$Q�E�$Q�E�$�MQ��$�UR�M��bE����tr�E$PQ�E �$Q�E�$Q�E�$�MQ�A�$�UR�M��/E����t?�E$PQ�E �$Q�E�$Q�E�$�MQ�A�$�UR�M���D����tǅ0���   �
ǅ0���    ��0���_^[���   ;������]�  �������������������������������������������������������������������U����   SVWQ��0����4   ������Y�M��E$PQ�E �$Q�E�$Q�E�$�MQ��$�UR�M��|@����tr�E$PQ�E �$Q�E�$Q�E�$�MQ�A�$�UR�M��I@����t?�E$PQ�E �$Q�E�$Q�E�$�MQ�A�$�UR�M��@����tǅ0���   �
ǅ0���    ��0���_^[���   ;��y����]�  �������������������������������������������������������������������U���  SVWQ�������B   ������Y�XD3ŉE��M�hCITb�M��:���EPhCITb�M��2���EPhsirt�M���B���EPhulav�M��B���E�P�MQ�����R�M��������-���������������'���M���
��������R��P��|����XZ_^[�M�3���/����  ;��[����]� �   �|����   �|msg ����������������������������������������������������������������������������U����   SVWQ������<   ������Y�M�j �EP�� ���Q�M���P�UR�M��A��������� ����	2�������_^[���   ;������]� ������������������������������U����   SVWQ��4����3   ������Y�M��EPj Q���$Q���$htemfQ�E�$Q�E�$Q�E�$Q�E�$�MQ�M��BC��_^[���   ;�������]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��EPj Q���$Q���$hrgdfQ�E�$��<���$Q�E�$��<���$Q�E�$��<���$Q�E�$�MQ�M��B��_^[���   ;��6����]� ������������������������������������������������U����   SVW��<����1   �������E�h.�5�Uٝ<���م<���_^[��]�����������������U����   SVWQ��(����6   ������Y�M��EPj Q���$Q���$htcpf�E�5�Uٝ0���م0���Q�$�E�5�Uٝ,���م,���Q�$�E�5�Uٝ(���م(���Q�$Q�E�$�MQ�M��\A��_^[���   ;������]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��I�M�l����P�EPQ�E�$Q�E�$�MQ�M�C;��P�U��BP��c�Q0�B4�Ѓ�;��W��_^[���   ;��G����]� �������������������������������������������������U����   SVWQ������9   ������Y�M��E��x u3��J�M�����P�E�P�M�:��P�M��QR��c�H0�Q8�҃�;�����E�3��}� ���M��E�R��P�������XZ_^[���   ;��u����]� �I    ������   ȁval ����������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��6�M�����P�EP�M�9��P�M��QR��c�H0�Q8�҃�;����_^[���   ;������]� ������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��6�M�����P�EP�M�9��P�M��QR��c�H0�Q<�҃�;����_^[���   ;��
����]� ������������������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M��t)����u3��;�E��P�MQ�M��Y)����u3�� �E��P�MQ�M��>)����u3���   _^[���   ;��Z����]� ������������������������������������U���   SVWQ�� ����@   ������Y�M��E��x u3��   �E�E�M������P�E�P�M�7��P�M��QR��c�H0�QD�҃�;������E��}� t\�}� tV�E�P�M��-���}� t=�E쉅������������������ tj������|���� ����
ǅ ���    �E�    �E�R��P������XZ_^[��   ;��8����]� ��   ������   �str ������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��*���E��t�E�P�b�����E�_^[���   ;��~����]� ������������������������U����   SVW��@����0   �������EP��c�Q�B�Ѓ�;��$��_^[���   ;������]���������������������������������U���  SVWQ�������C   ������Y�XD3ŉE��M�M������E�P�MQ�M��+���EЃ}� uǅ����    �M���(���������#�E�P�M�����EЉ�����M���(�������R��P������XZ_^[�M�3��%����  ;��:����]�    �����    �str ������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��;�M�|����P�EP�MQ�M�a4��P�U��BP��c�Q0�BH�Ѓ�;��u��_^[���   ;��e����]� �����������������������������������������������U����   SVWQ������9   ������Y�M��E�    �E�P�MQ�M��$���E��E�P�MQ�M����E�R��P�h��B��XZ_^[���   ;������]� �   p�����   |�b ��������������������������������������������������U����   SVWQ������9   ������Y�M��E�P�MQ�M�����E��E�P�MQ�M�%6���E�R��P� ����XZ_^[���   ;������]�    (�����   4�b ������������������������������������������U����   SVWQ������9   ������Y�M��E�P�MQ�M��T#���E�Q�E��$�EP�M�\����E�R��P�ԉ�� ��XZ_^[���   ;��S����]� �   ܉����   �b ��������������������������������������U����   SVWQ�� ����8   ������Y�M��M������E�P�MQ�M��"����u3��E�E�P�MQ�M��"����u3��-�E�P�MQ�M��l"����u3���E�P�MQ�M�A&���   R��P��������XZ_^[���   ;��g����]� �   Ȋ����   Ԋv ����������������������������������������������������������U���   SVWQ�� ����@   ������Y�XD3ŉE��M�M�����E�P�MQ�M��&���EЍE�P�MQ�M�x#���EЉ�����M��$�������R��P�������XZ_^[�M�3��� ����   ;��v����]�    ������   ċb ����������������������������������������������������������U���  SVWQ�������C   ������Y�XD3ŉE��M�M��|���E�P�MQ�M��*���EčE�P�MQ�M����Eĉ������M��T���������R��P�������XZ_^[�M�3��  ����  ;��
����]�    ������   ��b ����������������������������������������������������������U����   SVWQ������>   ������Y�M��M������E�P�M�Q�UR�M�������Ẽ}�t�E�P�MQ�M�#���}�tQ�E��$�EP�M�����E�R��P�������XZ_^[���   ;��	����]� �   ������   ������   ��b c ������������������������������������������������U����   SVWQ��4����3   ������Y�M�j j �EP�M���P�MQ�M�� ��_^[���   ;�������]� ��������������������������U����   SVWQ��4����3   ������Y�M��E$P�M Qj �UR�EP�MQj �UR�M�~1��P�EP�M�����_^[���   ;��l����]�  ��������������������������������������U����   SVWQ��4����3   ������Y�M�j �E,PQ�E(�$Q�E$�$�M QQ�E�$Q�E�$Q�E�$Q���$�UR�M� ��Q�$�EP�M��2��_^[���   ;������]�( ����������������������������������������U����   SVWQ��4����3   ������Y�M�j Q�E�$Q�E�$Q�E�$Q���$�EP�M�f��Q�$�MQ�M���(��_^[���   ;��$����]� ������������������������������U����   SVWQ��4����3   ������Y�M�j Q�E�$Q�E�$Q�E�$Q���$�EP�M����Q�$�MQ�M���.��_^[���   ;������]� ������������������������������U����   SVWQ��4����3   ������Y�M�j Q�E�$Q�E�$Q�E�$Q���$�EP�M�F��Q�$�MQ�M��*��_^[���   ;������]� ������������������������������U����   SVWQ������=   ������Y�M�j Q�E$�$Q�E �$Q�E�$��������P�EP��$���Q�M�,��P�UR�EP�MQ�M�����_^[���   ;��b����]�  ��������������������������������������������U����   SVWQ������=   ������Y�M�j Q�E$�$Q�E �$Q�E�$���������P�EP��$���Q�M�[+��P�UR�EP�MQ�M��(��_^[���   ;������]�  ��������������������������������������������U����   SVWQ������=   ������Y�M�j Q�E$�$Q�E �$Q�E�$������%��P�EP��$���Q�M�*��P�UR�EP�MQ�M����_^[���   ;������]�  ��������������������������������������������U����   SVWQ������=   ������Y�M�j Q�E$�$Q�E �$Q�E�$������u
��P�EP��$���Q�M��)��P�UR�EP�MQ�M������_^[���   ;��R����]�  ��������������������������������������������U���  SVWQ�������B   ������Y�M�j �EP������*��P�MQ�� ���R�M����P�EP�M���*���������� ����)����������������_^[��  ;������]� �����������������������������������U���   SVWQ�������H   ������Y�M�j ����������P�EP�����Q�M����P�UR�M��\���������������������������������_^[��   ;�������]� ���������������������������������������U���   SVWQ�� ����@   ������Y�M����]�}�tQ���$�EP�M�����]�EPQ�E�$Q�E��$������J��P�MQ�����R�M��'��P�EP�M��)��_^[��   ;��/����]� �����������������������������������������U���$  SVWQ�������I   ������Y�XD3ŉE��M�} u��c�H���   ��;�� ���E�} u3���  �M�����E�htlfv�M�����M�K%���M�ٝ����م����Q�$�=�����Mݝ�����$���Q�$�#����ܽ����ٝ����م����Q�$hulav�M�����hmrffhtmrf�M��(���M��$���M�ٝ����م����Q�$�������Mݝ��������Q�$�����ܽ����ٝ����م����Q�$hinim�M������M�y$���M�ٝ����م����Q�$�k�����Mݝ�����R���Q�$�Q����ܽ����ٝ����م����Q�$hixam�M��?���Q���$hpets�M��,���j hdauq�M��3'���E�Phspff�M��"'���E Phsirt�M��'���E�P�MQ������R�M��R����������������������C���M��5���������R��P�x��;���XZ_^[�M�3��(����$  ;�������]�    ������   ��msg ����������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��<����1   �������E���$������ٝ<���م<���_^[���   ;�������]����������������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U���  SVWQ�������B   ������Y�M��} u��c�H���   ��;������E�} u3��k�M������E�E�P�MQ�M��]���E��E���Nٝ����م����Q�$�E���Nٝ����م����Q�$������5�����P�E��P�E�R��P������XZ_^[��  ;��%�����]� �I    �����   �b ����������������������������������������������������������������������U����   SVWQ������;   ������Y�M�j �E P�MQ�UR��������P�EP��(���Q�M�c��P�UR�EP�M�����_^[���   ;��O�����]� �����������������������������������������U����   SVWQ������:   ������Y�M��M�����E�P�MQ�UR�M��N���E܍E�P�MQ�M�V����E�R��P�|��-���XZ_^[���   ;�������]�    ������   ��time �������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��D�M�������Pj j j j j j �M����Pj1�E��HQ��c�B0���   �у�(;������_^[���   ;��������]� ��������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj j �MQ�UR�EP�MQ�URj�E��HQ��c�B0���   �у�(;��7����E�R��P������XZ_^[���   ;�������]� �   �����   (�r ������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��7��j j j j j j j �EPj-�M��QR��c�H0���   �҃�(;��Y���_^[���   ;��I�����]� �����������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��F�E�    ��E�Pj j j �MQ�URj j j)�E��HQ��c�B0���   �у�(;������E�R��P�������XZ_^[���   ;�������]� �I    ������   ��r ����������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��F�E�    ��E�Pj j �MQj �URj j j)�E��HQ��c�B0���   �у�(;������E�R��P�������XZ_^[���   ;�������]� �I    ������   ��r ����������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��=��j j j �EP�MQ�URj �EPj/�M��QR��c�H0���   �҃�(;������_^[���   ;��������]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj j �MQ�UR�EP�MQ�URj'�E��HQ��c�B0���   �у�(;������E�R��P�4��v���XZ_^[���   ;��������]� �   <�����   H�r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj j �MQ�UR�EP�MQ�URj,�E��HQ��c�B0���   �у�(;��'����E�R��P�$�����XZ_^[���   ;�������]� �   ,�����   8�r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj j �MQ�UR�EP�MQ�URj�E��HQ��c�B0���   �у�(;��7����E�R��P������XZ_^[���   ;�������]� �   �����   (�r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��M�E�    ��E�Pj �MQ�UR�EP�MQ�UR�EPj�M��QR��c�H0���   �҃�(;��F����E�R��P������XZ_^[���   ;��"�����]�    �����   �r ������������������������������������������������������U����   SVWQ��4����3   ������Y�M���j j j �EP�MQ�URj �EPj.�M��QR��c�H0���   �҃�(;��p���_^[���   ;��`�����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj �MQ�UR�EP�MQj �URj�E��HQ��c�B0���   �у�(;������E�R��P�������XZ_^[���   ;�������]� �   ������   ��r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj �MQ�UR�EP�MQj �URj:�E��HQ��c�B0���   �у�(;�������E�R��P����&���XZ_^[���   ;�������]� �   ������   ��r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj �MQ�UR�EP�MQj �URj�E��HQ��c�B0���   �у�(;�������E�R��P�t��6���XZ_^[���   ;�������]� �   |�����   ��r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj �MQ�UR�EP�MQj �URj*�E��HQ��c�B0���   �у�(;�������E�R��P�d��F���XZ_^[���   ;��������]� �   l�����   x�r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��J�E�    ��E�Pj j �MQ�UR�EPj �MQj�U��BP��c�Q0���   �Ѓ�(;�������E�R��P�T��X���XZ_^[���   ;��������]� �I    \�����   h�r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��J�E�    ��E�Pj j �MQ�UR�EPj �MQj�U��BP��c�Q0���   �Ѓ�(;��	����E�R��P�D��h���XZ_^[���   ;��������]� �I    L�����   X�r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��J�E�    ��E�Pj j �MQ�UR�EPj �MQj	�U��BP��c�Q0���   �Ѓ�(;������E�R��P�4��x���XZ_^[���   ;��������]� �I    <�����   H�r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��J�E�    ��E�Pj j �MQ�UR�EPj �MQj
�U��BP��c�Q0���   �Ѓ�(;��)����E�R��P�$�����XZ_^[���   ;�������]� �I    ,�����   8�r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��J�E�    ��E�Pj j �MQ�UR�EPj �MQj�U��BP��c�Q0���   �Ѓ�(;��9����E�R��P������XZ_^[���   ;�������]� �I    �����   (�r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj �MQ�UR�EP�MQj �URj�E��HQ��c�B0���   �у�(;��G����E�R��P������XZ_^[���   ;��#�����]� �   �����   �r ������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��=��j j j �EP�MQ�URj �EPj�M��QR��c�H0���   �҃�(;��c���_^[���   ;��S�����]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj �MQ�UR�EP�MQj �URj�E��HQ��c�B0���   �у�(;������E�R��P�������XZ_^[���   ;�������]� �   ������   ��r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��J�E�    ��E�Pj j �MQ�UR�EPj �MQj�U��BP��c�Q0���   �Ѓ�(;������E�R��P�������XZ_^[���   ;�������]� �I    ������   ��r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��J�E�    ��E�Pj j �MQ�UR�EPj �MQj=�U��BP��c�Q0���   �Ѓ�(;�������E�R��P����(���XZ_^[���   ;�������]� �I    ������   ��r ������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��H�M�������Pj j j j �EP�MQ�M����Pj�U��BP��c�Q0���   �Ѓ�(;������_^[���   ;��������]� ��������������������������������������������������U����   SVWQ������=   ������Y�M��EP�M��>����E�P�M�Q�M��������t+�}� u��M��.���P�E�P�MQ�M�������u3�����   R��P�,�����XZ_^[���   ;��������]� ��   4�����   `�����   \�����   X�dat sid br �������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��D�M������Pj j j j j j �M����Pj�E��HQ��c�B0���   �у�(;�����_^[���   ;��������]� ��������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��J�E�    ��E�Pj j �MQ�UR�EPj �MQj�U��BP��c�Q0���   �Ѓ�(;��Y����E�R��P�������XZ_^[���   ;��5�����]� �I    ������   �r ������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��-��EP�MQ�UR�E��HQ��c�B0�HT�у�;�����_^[���   ;��s�����]� �����������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��9��EP�MQ�UR�EP�MQ�UR�E��HQ��c�B0�HX�у�;������_^[���   ;��������]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��!��E��HQ��c�B0�Hh�у�;��_���_^[���   ;��O�����]����������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��)��EP�MQ�U��BP��c�Q0�B\�Ѓ�;������_^[���   ;��������]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��)�E   ���P�M��QR��c�H0�Q`�҃�;��G���_^[���   ;��7�����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��$��EP�M��QR��c�H0�Q`�҃�;�����_^[���   ;�������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��0��EP�MQ�UR�EP�M��QR��c�H0�Qd�҃�;�� ���_^[���   ;�������]� ������������������������������������������U����   SVWQ��4����3   ������Y�M���E�HQ��c�B4��у�;������E�@    �E�M��H�M�V�����P�EP�MQ�M�;��P�U��BP��c�Q0���   �Ѓ�;��L����M�A�E3Ƀx ����_^[���   ;��(�����]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��7��j j j j j �EPj j j�M��QR��c�H0���   �҃�(;�����_^[���   ;��y�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��} u3��=�E�@    �M�7�����P�EP�M��(���P��c�Q0���   �Ѓ�;������_^[���   ;��������]� ��������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j0�M�����P��c�H0���   �҃�(;��V���_^[���   ;��F�����]�����������������������������������U����   SVWQ��4����3   ������Y�M��} u�E�c��EP�M�#���P�MQ�U��BP��c�Q0�BP�Ѓ�;�����_^[���   ;�������]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U��BP��c�Q0�Bt�Ѓ�;��(���_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U��BP��c�Q0���   �Ѓ�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M��M�	�����P�EP�MQ�UR�EP�M�����P�M��QR��c�H0�Qx�҃�;������_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j �M�Q���Pj�E��HQ��c�B0���   �у�(;��`���_^[���   ;��P�����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j jj �M����Pj�E��HQ��c�B0���   �у�(;������_^[���   ;�������]� ������������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j �M����Pj�E��HQ��c�B0���   �у�(;�� ���_^[���   ;�������]� ������������������������������������������U���  SVWQ�������A   ������Y�XD3ŉE��M�M��n����M�w�����P�E�Pj j j j j �M�V���Pj8�M�QR��c�H0���   �҃�(;��f����Ẽ}� t�E�P�M�m����Ẻ� ����M������� ���R��P������XZ_^[�M�3�������  ;�������]� �    �����   ,�storehere ��������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M�I�����P�EPj j j j j �M�(���Pj9�M��QR��c�H0���   �҃�(;��8���_^[���   ;��(�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��M������Pj j j j j j �M����Pj"�E��HQ��c�B0���   �у�(;�����_^[���   ;�������]� �����������������������������������U����   SVWQ��4����3   ������Y�M��M�	�����Pj j j j j j �M�����Pj5�E��HQ��c�B0���   �у�(;������_^[���   ;��������]� �����������������������������������U����   SVWQ��4����3   ������Y�M��M�i�����Pj j j j �EPj �M�H���Pj<�M��QR��c�H0���   �҃�(;��X���_^[���   ;��H�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���j j �EP�MQ�UR�EPj �MQj3�U��BP��c�Q0���   �Ѓ�(;�����_^[���   ;�������]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j �EPj �MQj�U��BP��c�Q0���   �Ѓ�(;��#�����EP�M��QR��c�H0���   �҃�;������_^[���   ;��������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j �EPj j�M��QR��c�H0���   �҃�(;��f���_^[���   ;��V�����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j�E��HQ��c�B0���   �у�(;������_^[���   ;��������]������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j �EPj�M��QR��c�H0���   �҃�(;��F���_^[���   ;��6�����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j(�E��HQ��c�B0���   �у�(;�����_^[���   ;�������]������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j �EP�MQj&�U��BP��c�Q0���   �Ѓ�(;��#���_^[���   ;�������]� �����������������������������U����   SVWQ��4����3   ������Y�M���j j j j �EP�MQj �URj+�E��HQ��c�B0���   �у�(;�����_^[���   ;�������]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j�E��HQ��c�B0���   �у�(;������_^[���   ;��������]������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j#�E��HQ��c�B0���   �у�(;��g���_^[���   ;��W�����]������������������������������������U����   SVWQ��4����3   ������Y�M��} tj j�M������M��} tj j�M������M���EP�MQ�U��BP��c�Q0�Bp�Ѓ�;�����_^[���   ;�������]� ������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E��HQ��c�B0���   �у�;�����_^[���   ;�������]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j �E��HQ��c�B0���   �у�(;�����_^[���   ;��w�����]������������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]������������������U����   SVWQ��4����3   ������Y�M��   _^[��]������������������U����   SVWQ��4����3   ������Y�M�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M��M������E�� �U�E��@   �E��@    �E�_^[���   ;��5�����]����������������������������������U����   SVWQ��4����3   ������Y�M��M��H����E��t�E�P�m������E�_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� �U�M��r���_^[���   ;��\�����]�������������������������U����   SVWQ��0����4   ������Y�M�j �EP�MQ�UR�EPj j �M�������t�M��y tǅ0���   �
ǅ0���    ��0���_^[���   ;��������]� ��������������������������������U����   SVWQ��4����3   ������Y�M��E��M�H�M��	���_^[���   ;��\�����]� ����������������������U����   SVWQ������:   ������Y�M��M��������������ckhc)�����ckhct5�����cksatY�����TCAbtr��   �����atnit��   3���   �E��x t �M�������t�E��@    �   �   3��   �E��x t�E����M��B��;��s����}3��yj hdiem�M�S����E�E��@   ��EP�M�Q�U���M��P��;��3����E��E��x t�}�t�}�u3��}���P�M������E���EP�MQ�M��ν��_^[���   ;��������]� ����������������������������������������������������������������������������������������������U����   SVWQ�� ����8   ������Y�M��E��x u�  �E�� ����� �����   �� ����$����E;E~��   �   �E;E|��   �{�E;E}�   �l�E;E�   �]�E;E~�E;E}�   �F�E;E|
�E;E�x�2�E;E|
�E;E}�d��E;E~
�E;E�P�
�E;Et�D�EP��(����w�����(���Q�M�����j�EQ�$�EQ�$�EP�������E��@    _^[���   ;��<�����]� ������$�3�J�^�r���������������������������������������������������������������������������������������������������U����   SVWQ�� ����8   ������Y�M��E��x u�l  �E�� ����� ����  �� ����$�$��E�E������z�5  ��   �E�E������Az�  ��   �E�E������Au�  �   �E�E������u��   �   �E�E������z�E�E������Au��   �z�E�E������Az�E�E������u�   �U�E�E������Az�E�E������Au�{�3�E�E������z�E�E������u�Y��E�E������D{�F�EP��(����@�����(���Q�M��o����EPQ�E�$Q�E�$�MQ�ټ�����E��@    _^[���   ;�������]� ��������(�M�r�����������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�jQ�E�$Q�E�$Q�E�$�EP�MQ�M��1���_^[���   ;�������]� ��������������������������������U����   SVWQ��4����3   ������Y�M�jQ�E�$Q�E�$Q�E�$�EP�MQ�M�豳��_^[���   ;�膿����]� ��������������������������������U����   SVWQ��4����3   ������Y�M�jQ�E�$Q�E�$Q�E�$�EP�MQ�M��1���_^[���   ;�������]� ��������������������������������U����   SVWQ��4����3   ������Y�M��E�� �U�E��@    �E��@    �E��@    �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��M��P����E��t�E�P�ͱ�����E�_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� �U�E��x u ��E��HQ��c�B4��у�;�諽���E��@    �E��@    _^[���   ;�臽����]������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��c�H4�Qx�҃�;�����_^[���   ;��	�����]� �����������������������������������U����   SVWQ��(����6   ������Y�M��} tT��EP�M��Ϲ��P��c�Q0���   �Ѓ�;�荼���E��EP�M�Q��c�B0���   �у�;��e����'��EP�M��QR��c�H0���   �҃�;��<���_^[���   ;��,�����]� ������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��c�B4�H�у�;�謻��_^[���   ;�蜻����]�������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��c�B4�H�у�;��<���_^[���   ;��,�����]�������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��c�B4�H�у�;��̺��_^[���   ;�輺����]�������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��c�B4���   �у�;��Y���_^[���   ;��I�����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��c�B4���   �у�;��ٹ��_^[���   ;��ɹ����]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��QR��c�H4�Q�҃�;��M���_^[���   ;��=�����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��QR��c�H4�Q�҃�;�轸��_^[���   ;�譸����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��c�H4�Q �҃�;��9���_^[���   ;��)�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��c�H4�Q$�҃�;�蹷��_^[���   ;�詷����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��QR��c�H0���   �҃�;��*���_^[���   ;�������]� ������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��c�H4���   �҃�;�覶��_^[���   ;�薶����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U��BP��c�Q4���   �Ѓ�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U��BP��c�Q4���   �Ѓ�;�腵��_^[���   ;��u�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��c�H4�Q(�҃�;��	���_^[���   ;��������]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E��HQ��c�B4�H,�у�;�耴��_^[���   ;��p�����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��c�Q4�B0�Ѓ�;�����_^[���   ;��������]� ������������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��c�B4�H4�у�;�茳��_^[���   ;��|�����]�������������������������U���(  SVWQ�������J   ������Y�M��E�    �E�    �E�P�M�Q�UR�E��H�����M�����P������������E�P�M�Q�U�R�E�P������Q�U��J������} tL�} tF�E�;E�~*�M�M�9M�}�U�;U�~�E�E�9E�}ǅ����   �
ǅ����    �������h�7�} t1�E�;E�~�M�M�9M�}ǅ����   �
ǅ����    �������/�E�;E�~�M�M�9M�}ǅ����   �
ǅ����    ������R��P� �茥��XZ_^[��(  ;��	�����]� �I    (�����   |�����   z�����   x�����   v�����   s�����   p�dy dx h w y x ������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��c�H4�Q8�҃�;�����_^[���   ;��ٰ����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��c�H4�Q<�҃�;��i���_^[���   ;��Y�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��c�Q4���   �Ѓ�;�����_^[���   ;��ѯ����]� ���������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��c�B4�H@�у�;��l���_^[���   ;��\�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��c�Q4�BD�Ѓ�;������_^[���   ;�������]� ������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��c�Q4�BH�Ѓ�;��t���_^[���   ;��d�����]� ������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��c�Q4�BL�Ѓ�;������_^[���   ;�������]� ������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��c�Q4�BP�Ѓ�;��t���_^[���   ;��d�����]� ������������������������������U����   SVWQ��4����3   ������Y�M��M耺����u�-��EP�MQ�UR�E��HQ��c�B4�HT�у�;�����_^[���   ;��Ҭ����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M���E,P�M(Q�U$R�E P�MQ�UR�EP�MQ�UR�EP�M��QR��c�H4�QX�҃�,;��5���_^[���   ;��%�����]�( �����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��QR��c�H4�Q\�҃�;�蝫��_^[���   ;�荫����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��c�B4�Hd�у�;�����_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��c�B4�Hh�у�;�謪��_^[���   ;�蜪����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR�E��HQ��c�B4�H`�у�;��$���_^[���   ;�������]� ������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��c�Q4�Bl�Ѓ�;�褩��_^[���   ;�蔩����]� ������������������������������U����   SVWQ��(����6   ������Y�M��} t�E��ًU�
�} t�E��ًU�
��EP�MQ�U��BP��c�Q4�Bl�Ѓ�;�� ����E�} t�E��ًU�
�} t�E��ًU�
�E�_^[���   ;��ƨ����]� ������������������������������������������������U����   SVWQ��(����6   ������Y�M��} t�E��ًU�
�} t�E��ًU�
��EP�MQ�U��BP��c�Q4�Bt�Ѓ�;�� ����E�} t�E��ًU�
�} t�E��ًU�
�E�_^[���   ;�������]� ������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��c�Q4�Bt�Ѓ�;��d���_^[���   ;��T�����]� ������������������������������U���  SVWQ�������B   ������Y�M��E��x ��   �} t4�M�衻����P�E��H�
���P��c�Q0���   �Ѓ�;��Ȧ���T�M��m���P�����訦��hARDb����������P�����P��(���Q�U��J�ۙ����(����ٳ���������Ȗ��_^[��  ;��b�����]� ������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��c�H4�Qp�҃�;��٥���   _^[���   ;��ĥ����]� ������������������������������U����   SVWQ��4����3   ������Y�M���EPQ�E�$Q�E�$�MQ�U��BP��c�Q4���   �Ѓ�;��C���_^[���   ;��3�����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E��HQ��c�B4���   �у�;�轤��_^[���   ;�譤����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��c�B4���   �у�;��9���_^[���   ;��)�����]��������������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]������������������U����   SVWQ��4����3   ������Y�M��   _^[��]������������������U����   SVWQ��4����3   ������Y�M�h�  �M��!����EP�MQ�UR�EP�M�����2�_^[���   ;��&�����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M���M��B��;�跢��_^[���   ;�觢����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��QR��c�H4�Q|�҃�;�����_^[���   ;��ݠ����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�UR�E��H�ò��_^[���   ;��f�����]� ��������������������������������U����   SVWQ��4����3   ������Y�M��} tj j�M� ����M��} tj j�M������M���EP�MQ�U��BP��c�Q4�Bt�Ѓ�;��Ɵ��_^[���   ;�趟����]� ������������������������������������������������U���0  SVWQ�������L   ������Y�M��E�    �M����������������INIbf������INIb��   ������SACb5������SACb��   ������$'  ��  ������MicM��  �$  ������ARDb�4  �  ������NIVb1������NIVbt\������NPIb�v  ������ISIb��   ��  ������cnys��  �  �E����M��B��;��n����E�   �  �E����M��B��;��L����E�   �y  �E�    �E�    ��E�P�M�Q�U���M��P��;�������t)��E�P�M�Q�U��BP��c�Q4�B�Ѓ�;������E�   �  �M��d�����P�M�轔��P�E���M��B��;�賝���E�   ��   j j�M�����E�j j�M�����E�j j�M�r����E�j j�M�c����E���EP�M�Q�U�R�E�P�M�Q�U���M��P��;��A����E�   �q��EP�M���M��B��;������X��EP�M���M��B$��;������E�   �2j hIicM�M������E��EP�M�Q�U���M��P ��;��ɜ����E�R��P����&���XZ_^[��0  ;�補����]� �   ������   ������   ��h w ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�h����h����h�����EP�MQh����h����h����h�����UR�M��{���_^[���   ;��F�����]� ��������������������������������U����   SVWQ������:   ������Y�M�hYALf����������P�M��|���������/���_^[���   ;��ɚ����]��������������������������������������U����   SVWQ��4����3   ������Y�M��M��ě���E�� 4V�E��@   �E�_^[���   ;��O�����]����������������������������U����   SVWQ��4����3   ������Y�M��M�舞���E��t�E�P荍�����E�_^[���   ;��ޙ����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� 4V�M�蒘��_^[���   ;��|�����]�������������������������U����   SVWQ��0����4   ������Y�M��M�ڷ����0�����0���cksat9��0���ckhct�P�E��@   �M��S�����t�E��@    �   �93��5�E��x t�E����M��B��;��˘���3���EP�MQ�M�菑��_^[���   ;�襘����]� ���������������������������������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR��c�H��H  �҃�;�����_^[���   ;��������]���������������������������U����   SVW��@����0   �������EP��c�Q0���   �Ѓ�;�街��_^[���   ;�著����]������������������������������U����   SVW��(����6   �������EP�MQ��,���R��c�H0���   �҃�;��'���P�M� �����,���肯���E_^[���   ;�� �����]���������������������������������������������U���0  SVW�������L   ������XD3ŉE��M��ޞ���E�    �	�E܃��Eܸ   ����   j �E�k�
P�M�e����E�j �E�k�
��P�M�N����Eă}� u�b�}� ~,j h`V�������4���������P�M��H���������苮���E�P�M�Q������R������P�M������������`����U����E�P�M�����M��G����ER��P�|�7���XZ_^[�M�3��$�����0  ;�誕����]Ë�   �����   �t ����������������������������������������������������������������������������������������������U����   SVW��@����0   �������EP�MQ��c�B0���   �у�;�����_^[���   ;��ݔ����]��������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR��c�H0���   �҃�;��n���_^[���   ;��^�����]���������������������������U����   SVW��@����0   ������j0�EP�̱����_^[���   ;�������]�����������������U����   SVW��@����0   ������j0�EP������P�s�����_^[���   ;�諓����]������������������������U����   SVW��(����6   ������j0�EP�MQ��,���R�&�����P��������,���贫��_^[���   ;��5�����]����������������������������������U����   SVW��(����6   ������j0�EP�MQ�UR��,���P�_�����P脰������,����0���_^[���   ;�豒����]������������������������������U����   SVW��@����0   ������j$�EP������3Ƀ�����_^[���   ;��J�����]�����������������������U����   SVW��@����0   ������j$�EP�Q����P賯����3Ƀ�����_^[���   ;�������]������������������������������U����   SVW������9   ������j$�EP�MQ��,���R�V�����P�8�����3Ƀ����� �����,����֩���� ���_^[���   ;��Q�����]������������������������������U����   SVW������9   ������j$�EP�MQ�UR��,���P������P褮����3Ƀ����� �����,����B����� ���_^[���   ;�轐����]������������������������������������������U����   SVW��@����0   �������EP�MQj ��c�B��  �у�;��K���_^[���   ;��;�����]������������������������U����   SVW��@����0   �������EP�MQ�URj ��c�H��  �҃�;��؏��_^[���   ;��ȏ����]�������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E��HQ��c�B4�H,�у�;��P���_^[���   ;��@�����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��c�Q4�B0�Ѓ�;��Ԏ��_^[���   ;��Ď����]� ������������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��c�B4�H4�у�;��\���_^[���   ;��L�����]�������������������������U����   SVWQ������9   ������Y�M��M��~��� �E�M�`����E��}� t�E�   �E�P�M�Q�UR�M��n���_^[���   ;��č����]� ������������������������������U����   SVWQ��4����3   ������Y�M��E P�MQ�M�N���P�UR�EP�MQ�M�֑���R�EP�M�賖��_^[���   ;��9�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��M�;x��P�E(PQ�E$�$Q�E �$�MQQ�E�$Q�E�$Q�E�$�M�3���Q� �$�UR�M�����_^[���   ;�菌����]�$ �����������������������������������������U����   SVWQ��4����3   ������Y�M��M�w��PQ�E�$Q�E�$Q�E�$�M虯��Q� �$�EP�M�豭��_^[���   ;��������]� �������������������������������U����   SVWQ��4����3   ������Y�M��M��v��PQ�E�$Q�E�$Q�E�$�M�	���Q� �$�EP�M�蘳��_^[���   ;��e�����]� �������������������������������U����   SVWQ��4����3   ������Y�M��M�kv��PQ�E�$Q�E�$Q�E�$�M�y���Q� �$�EP�M��R���_^[���   ;��Պ����]� �������������������������������U����   SVWQ��4����3   ������Y�M��M茦��P�EP�MQ�UR�M芬��P�EP�MQ�M�����_^[���   ;��O�����]� �������������������������U����   SVWQ��4����3   ������Y�M��M�\���PQ�E �$Q�E�$Q�E�$�M�z���P�EP�MQ�UR�M��8���_^[���   ;������]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M輠��PQ�E �$Q�E�$Q�E�$�M�ڠ��P�EP�MQ�UR�M�蘌��_^[���   ;��"�����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M����PQ�E �$Q�E�$Q�E�$�M�:���P�EP�MQ�UR�M��&���_^[���   ;�肈����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M�|���PQ�E �$Q�E�$Q�E�$�M蚟��P�EP�MQ�UR�M��cq��_^[���   ;�������]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M����P�M����P�MQ�M��u���_^[���   ;��[�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��EPQ�E�$Q�E�$�M膞��P�MQ�M��В��_^[���   ;��ֆ����]� ��������������������������������U���  SVWQ�������F   ������Y�M��E�P�M�Q�UR�M������E�P�M�Q�U�R�E�P�MQ�M��c����} tL�} tF�E�;E�~*�M�M�9M�}�U�;U�~�E�E�9E�}ǅ����   �
ǅ����    �������h�7�} t1�E�;E�~�M�M�9M�}ǅ����   �
ǅ����    �������/�E�;E�~�M�M�9M�}ǅ����   �
ǅ����    ������R��P���y��XZ_^[��  ;�脅����]� ��   �����    ����   �����   �����   �����   �����   �dy dx h w y x ��������������������������������������������������������������������������������������������������������������U����   SVWQ������9   ������Y�M��E�E�}� u	�E����E�j hdiuM�M�^����E��}� u�   �G�E�M�;u3��9j hIicM�M�1���9E�uj h1icM�M������t3���E�M���   _^[���   ;�������]� ������������������������������������������������������������U����   SVW������:   ������hfnic�M�@~���E��}� tj
�M�蕄�����t�\hfnic�����P�M�u��P�M�z���������s���M�������t�M������uhfnic�M�ڣ���EPj
�M�ߚ��_^[���   ;�������]������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M����P��c�Q0���   �Ѓ�;��w���_^[���   ;��g�����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j6�M��'��P��c�H0���   �҃�(;�����_^[���   ;��ց����]�����������������������������������U����   SVWQ��(����6   ������Y�M�j �EP�M�~���E�E�P�M��en��_^[���   ;��`�����]� ��������������������������U����   SVWQ��(����6   ������Y�M�j �EP�M�����E�E�P�M�����_^[���   ;��������]� ��������������������������U����   SVWQ��(����6   ������Y�M�Q���$�EP�M�|���]�Q�E��$�M��ؚ��_^[���   ;��y�����]� �����������������������������������U���  SVWQ�������B   ������Y�M��M���������������P�EP�����Q�M芦����U�H�M�P�U���ċM��U�P�M�H�M��cv��R��P�p�9s��XZ_^[��  ;������]�    x����   �val ��������������������������������������������������������U����   SVWQ������?   ������Y�M��M��B���������7���P�EP�����Q�M�	�����@�U�E�E�P�M�Q�M��}��R��P�L�]r��XZ_^[���   ;���~����]�    T����   `val ��������������������������������������������U���$  SVWQ�������I   ������Y�XD3ŉE��M�M�虆��������莆��P�EP������Q�M�7���P�M��r���������藖��������茖�����̍E�P�����M��o���M��n���R��P�T�aq��XZ_^[�M�3��N�����$  ;���}����]� ��   \����   hval ��������������������������������������������������������������������U����   SVWQ������:   ������Y�M��E;Eu&j htsem�M�+�����uj hrdem�M������t3��B�E�    �EP�������|���M�Q�����R�M�
�����u3���E�P�M���i���   R��P�p�;p��XZ_^[���   ;��|����]� ��   x����   �val ��������������������������������������������������������U����   SVWQ������:   ������Y�M��E;Eu&j htsem�M������uj hrdem�M������t3��B�E�    �EP�������{���M�Q�����R�M�Z|����u3���E�P�M���}���   R��P���+o��XZ_^[���   ;��{����]� ��   �����   �val ��������������������������������������������������������U����   SVWQ������:   ������Y�M��E;Eu&j htsem�M������uj hrdem�M�������t3��C���]�EP�������z���M�Q�����R�M蛐����u3��Q�E��$�M������   R��P���n��XZ_^[���   ;��z����]� �   �����   �val ��������������������������������������������������������U���  SVWQ�������D   ������Y�M��E;Et�E;Et�E;Et3��   j htsem�M������uj hrdem�M�Ѣ����t3��   Q���$�M��W|���EP�������y���MQ������y���UR������y���E�P������Q�����R�����P�M�a�����u3��#���ċM��U�P�M�H�M���o���   R��P� �l��XZ_^[��  ;��)y����]� �I    ����   val ����������������������������������������������������������������������������������������U����   SVWQ������;   ������Y�M��E;Eu&j htsem�M�k�����uj hrdem�M�X�����t3��K�M��`���EP������:x���M�Q�UR�����P�M蚒����u3���E�P�M�Q�M���v���   R��P�8�rk��XZ_^[���   ;���w����]� �   @����   Lval ����������������������������������������������������������������U���  SVWQ�������G   ������Y�XD3ŉE��M�E;Eu&j htsem�M�A�����uj hrdem�M�.�����t3��v�M��g���EP�������w���M�Q������R�M������uǅ����    �M��`����������.���̍E�P�݃���M��;x��ǅ���   �M��0��������R��P�� �j��XZ_^[�M�3��
�����  ;��v����]� ��   � ����   � val ��������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��6����E�� lV�E��M�Hj hmyal�M�ɞ���M��A�E��xt�E��xt
�E��@    j hhfed�M蘞���M��A�E�_^[���   ;��u����]� ����������������������������������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�h�����E�_^[���   ;���t����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��8y��_^[���   ;��t����]������������������U����   SVWQ��0����4   ������Y�M��M�
�����0�����0���ytsdt�%�M��҆���E����M��B��;��3t���   ��EP�MQ�M���{��_^[���   ;��t����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ�� ����8   ������Y�M��M��f`���E�P�M�����M�諉���ER��P�l%�@e��XZ_^[���   ;��q����]� �I    t%����   �%tri ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M����~��_^[���   ;��2q����]�������������������������������U����   SVWQ��4����3   ������Y�M��E��M���E��P�M����Dq���E�_^[���   ;��p����]� ������������������������U����   SVWQ��4����3   ������Y�M��E����M��BD��;��gp����t*�E��H;Mt�E��M�H�E����M��BH��;��9p��_^[���   ;��)p����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��x u3���E��H��������_^[��]�������������������������U����   SVWQ��4����3   ������Y�M�_^[��]�����������������������U����   SVWQ��$����7   ������Y�M��M����[���E�� ������(����[��P�M����c[����(����#|���E�_^[���   ;��n����]���������������������������������U����   SVWQ��4����3   ������Y�M��E�3Ƀ8����_^[��]��������������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��8�u�E��     �E��M�H��E��8 u�E��H;Mt	�E��    _^[��]� ����������������������������U����   SVWQ��4����3   ������Y�M��E�3Ƀ8����_^[��]��������������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��(����6   ������Y�M��E��8�u�E��     �EP�M��������$�E��8 u�EP�M����8n����t	�E��    �M����R��P��*��_��XZ_^[���   ;��^l����]�    �*����   �*_$ArrayPad ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E�3Ƀ8����_^[��]��������������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��8�u�E��     �E��M�H��E��8 u�E��H;Mt	�E��    _^[��]� ����������������������������U����   SVWQ��4����3   ������Y�M��E�3Ƀ8����_^[��]��������������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��8�u�E��     �E��E�X�#�E��8 u�E��@�E������D{	�E��    _^[��]� �������������������������������������U����   SVWQ��4����3   ������Y�M��E�3Ƀ8����_^[��]��������������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��8�u"�E��     �E����M��U�P�M�H�(�E��8 u �EP�M���Q��f������t	�E��    _^[���   ;��h����]� �������������������������������������U����   SVW��<����1   ������E� �M�������Dz6�U�B�E�@������Dz!�M�A�U�B������Dzǅ<���    �
ǅ<���   ��<���_^[��]�����������������������������������U����   SVWQ��4����3   ������Y�M��E�3Ƀ8����_^[��]��������������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��8�u�E��     �E��M�H�U�P�(�E��8 u �EP�M���Q�P������t	�E��    _^[���   ;���f����]� ���������������������������������������������U����   SVW��,����5   ������E� �M�������Dz�E�@�M�A������Dz3��w�E� �M�Iٝ<���م<���Q�$�|�����U��E�Hٝ8���م8���Q�$ݝ0�����{����݅0���������D{ǅ,���   �
ǅ,���    ��,���_^[���   ;���e����]������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M������_^[��]� ���������������U����   SVWQ��4����3   ������Y�M������_^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��E�     _^[��]� ���������������������������U���  SVW��x����b   ������} u3��vj h�   ��<���P�i����ǅ@������E��<����E��\���ǅ|���3��E�0��E����E���E�ݢh�   ��<���P�MQ�URj轂����R��P��4�V��XZ_^[�Ĉ  ;��b����]Ð   �4<����   �4np ���������������������������������������������������������������������U���  SVW��x����b   ������} u3��   j h�   ��<���P�h����ǅ@������E��<����E��\����E��|����E�3��E����E�0��E���E�ݢ�E�{�h�   ��<���P�MQ�URj荁����R��P��5��T��XZ_^[�Ĉ  ;��aa����]Ð   �5<����   �5np ���������������������������������������������������������������������U����  SVW������z   ������M�En����tj �EP�MQ�L������u3��dj h   ������P�Rg�����EPj j �MQ�UR������P� m����ǅ|������E���h   ������P�MQ�URj�c�����R��P��6�S��XZ_^[���  ;��7`����]ÍI    �6����   7np ���������������������������������������������������������U����  SVW������z   ������M�%m����tj �EP�MQ�K������u3��cj h   ������P�2f�����E Pj j �MQ�UR������P��k�����E��|����E���h   ������P�MQ�URj�D����R��P�8�R��XZ_^[���  ;��_����]�   8����    8np ������������������������������������������������������������̋�`����������̋�`@����������̋�`����������̋�`����������̋�`D����������̋�`����������̋�`����������̋�`�����������U����   SVWQ��4����3   ������Y�M��E��@    �M��    �E��@    �E��@   �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��} u�4�} t�EP�M�t��� �} t�EP�M�LO����E�P�M�>O��_^[���   ;��a]����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP��c���   �M��B@��;���\��_^[���   ;���\����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��c���   �M��BD��;��|\��_^[���   ;��l\����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��c�Q@�M����   ��;��\��_^[���   ;���[����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��c�Q@�M����   ��;��[��_^[���   ;��[����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��c�B@�M����   ��;��([��_^[���   ;��[����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��c�B@�M����   ��;��Z��_^[���   ;��Z����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP��c���   �M����   ��;��)Z��_^[���   ;��Z����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��c���   �M����   ��;��Y��_^[���   ;��Y����]� �������������������������������U����   SVWQ��4����3   ������Y�M���c�P@��M����   ��;��1Y��_^[���   ;��!Y����]������������������������������U����   SVWQ��4����3   ������Y�M���c�P@��M����   ��;���X��_^[���   ;��X����]������������������������������U����   SVWQ��4����3   ������Y�M���EP��c�Q@�M����   ��;��LX��_^[���   ;��<X����]� ����������������������U����   SVWQ��4����3   ������Y�M���c�P@��M����   ��;���W��_^[���   ;���W����]������������������������������U����   SVWQ��4����3   ������Y�M���c���   ��M��Bt��;��qW��_^[���   ;��aW����]������������������������������U����   SVWQ��4����3   ������Y�M���EP��c�Q@�M����   ��;���V��_^[���   ;���V����]� ����������������������U����   SVWQ��(����6   ������Y�M���E�P��c�Q@�B$�Ѓ�;��V���E�E�#Et�E��#E�E��	�E�E�E��E�P�M�Q��c�B@�H �у�;��LV��_^[���   ;��<V����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH���   �Ѓ�;���U��_^[���   ;��U����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B@���   �у�;��XU��_^[���   ;��HU����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q@���   �Ѓ�;���T��_^[���   ;���T����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q@�B,�Ѓ�;��oT��_^[���   ;��_T����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B@�H(�у�;���S��_^[���   ;���S����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q@�BP�Ѓ�;��sS��_^[���   ;��cS����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B@�HT�у�;���R��_^[���   ;���R����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H@�QX�҃�;��xR��_^[���   ;��hR����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B@�H\�у�;���Q��_^[���   ;���Q����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��c���   �M��P��;��xQ��_^[���   ;��hQ����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��c���   �M��B��;���P��_^[���   ;���P����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��c���   �M��B ��;��uP��_^[���   ;��eP����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP��c���   �M����   ��;���O��_^[���   ;���O����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQQ�E�$�UR�EP�MQ��c���   �M����   ��;��RO��_^[���   ;��BO����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ��c���   �M����   ��;��N��_^[���   ;��N����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���c���   ��M��B$��;��AN��_^[���   ;��1N����]������������������������������U����   SVW��@����0   �����󫡨c�H@��Ql��;���M��_^[���   ;���M����]�������������������������U����   SVW��@����0   �������j�EPj ��c�Q@�Bp�Ѓ�;��pM��_^[���   ;��`M����]�����������������������������U����   SVW��@����0   �������j�EPh   @��c�Q@�Bp�Ѓ�;���L��_^[���   ;���L����]��������������������������U����   SVW��@����0   �������EP�MQj ��c�B@�Hp�у�;��L��_^[���   ;��~L����]���������������������������U����   SVW��@����0   �����󫡨c���   ����;��*L��_^[���   ;��L����]�����������������������U����   SVW��@����0   ������E�8 t#��E�Q��c���   �H�у�;��K���E�     _^[���   ;��K����]���������������������������U����   SVW��@����0   �����󫡨c���   ��Q ��;��IK��_^[���   ;��9K����]����������������������U����   SVW��@����0   ������E�8 t#��E�Q��c���   �H(�у�;���J���E�     _^[���   ;��J����]���������������������������U����   SVW��@����0   �����󫡨c�H@��Ql��;��lJ��_^[���   ;��\J����]�������������������������U����   SVW��@����0   ������E�8 t ��E�Q��c�B@�HH�у�;���I���E�     _^[���   ;���I����]������������������������������U����   SVW��@����0   �������EP��c�Q@���   �Ѓ�;��I��_^[���   ;��qI����]������������������������������U����   SVW��@����0   ������E�8 t ��E�Q��c�B@�HH�у�;��
I���E�     _^[���   ;���H����]������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QH���   �Ѓ�;��H��_^[���   ;��|H����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BH���  �у�;��H��_^[���   ;��H����]� ����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��c�Q �Bd�Ѓ�;��G��_^[���   ;��G����]�������������������������������������U����   SVW��4����3   ������}qF t�1�E�E��}� u�#�EP�M���8���E�P�MQ�M�c������[��_^[���   ;���F����]�����������������������������������U����   SVWQ��4����3   ������Y�M���c�P@��M����   ��;��F��_^[���   ;��F����]������������������������������U����   SVWQ��4����3   ������Y�M���EP��c�Q@�M����   ��;��F��_^[���   ;��F����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��c�B@�M����   ��;��E��_^[���   ;��E����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���c�P@��M����   ��;��1E��_^[���   ;��!E����]������������������������������U���(  SVWQ�������J   ������Y�M��E�� ��.����z�M����ٝ������U��ٝ����م�����]�E��@��.����z�M��A��ٝ������U��Bٝ����م�����]��E��8O����{�E��8O����z�E�����E����X�>  �E���V����zc�E���V����zS�E��f���E��E��f���E��Eș�}��U��E��EȋE��E��}� u��EȋE��8�M���EȋE��x�M��Y��   �E����$�E���$�aD�����=�V�]����]�����Au.�E��M��]��E��M��]��E�� �M��M���E��@�M��M��Y�E��X.����z���]��E����XQ�E��$Q�E��$�Q�����]��E��]��E��]��E���N����tˋE�� �u�M���E��@�u�M��Y_^[��(  ;���B����]�������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �������E�]����Au�E��E_^[��]�����������������������U����   SVW��<����1   �������E���$�E���$��P����ٝ<���م<���_^[���   ;��A����]�������������������������U����   SVW��@����0   �������EP��c�Q ���   �Ѓ�;��aA��_^[���   ;��QA����]������������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;���@���E�     _^[���   ;���@����]��������������������������������������U����   SVW��@����0   �����󫡨c�H ����;��}@��_^[���   ;��m@����]��������������������������U����   SVW��@����0   ������E�8 u�)��E�Q��c�B �H�у�;��@���E�     _^[���   ;���?����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B �HP�у�;��?��_^[���   ;��{?����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B �H�у�;��?��_^[���   ;���>����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B �H�у�;��>��_^[���   ;��{>����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q �B�Ѓ�;��>��_^[���   ;���=����]����������������������������U����   SVWQ������;   ������Y�XD3ŉE��M�M��n*����E�P�M�Q��c�B �H �у�;��=���E�P�M�g���M���-���ER��P��Y��0��XZ_^[�M�3���R�����   ;��G=����]� �   �Y����   �Ybc ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B �H$�у�;��<��_^[���   ;��<����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q �BD�Ѓ�;��/<��_^[���   ;��<����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q �BL�Ѓ�;��;��_^[���   ;��;����]����������������������������U����   SVWQ��4����3   ������Y�M��M��t'���E�� �V�E��@    �E�_^[���   ;��?;����]����������������������������U����   SVWQ��4����3   ������Y�M��M��_S���E��t�E�P�}.�����E�_^[���   ;���:����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��4��_^[���   ;��u:����]������������������U����   SVWQ��4����3   ������Y�M��E��M�H�   _^[��]� ����������������������U����   SVWQ��4����3   ������Y�M��E��x tj�EP�M��I�?���EP�MQ�M���O��_^[���   ;��9����]� �����������������������������U����   SVWQ��4����3   ������Y�M��E� P   �M�P   �   _^[��]� �����������������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M��M�����6���E��     �E��@    �E��@    �E�_^[���   ;��8����]�������������������������������U����   SVWQ��4����3   ������Y�M��E��8 t ��E��Q��c�B �H4�у�;��%8���M����P��_^[���   ;��
8����]���������������������������������������U����   SVWQ��$����7   ������Y�M��E��M�H�M��4���M��A�E��x u3��   �E�P�M����O$���}( t'�E(P��(����h7��j��(���Q�U���R�M�4N����E0P�M,Q�U(R�E$P�M Q�UR�EP�MQ�UR�M����)(��P�M�F4��P�E��HQ��c�B �H0�у�0;�� 7���U���E�3Ƀ8 ����_^[���   ;���6����]�, ������������������������������������������������������������������������U����   SVWQ������;   ������Y�XD3ŉE��M�E�8 u�B�M��#��hNIVb�M���V����j �E�P�M�R��c�H �Q8�҃�;��6���M��m&��R��P�8a�y)��XZ_^[�M�3��fK�����   ;���5����]�   @a����   Lamsg ������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 t�E��x t	�E��x u3��(��EP�MQ�U��P��c�Q �B8�Ѓ�;��75��_^[���   ;��'5����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QD�B�Ѓ�;��4��_^[���   ;��4����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QD�B�Ѓ�;��O4��_^[���   ;��?4����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QD�BP�Ѓ�;���3��_^[���   ;���3����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QD�B�Ѓ�;��o3��_^[���   ;��_3����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QD�B(�Ѓ�;���2��_^[���   ;���2����]����������������������������U����   SVWQ�� ����8   ������Y�M���E�P��$���Q��c�BX��у�;��2���U��
�H�J�@�B�E_^[���   ;��c2����]� �����������������������������U����   SVWQ�� ����8   ������Y�M���E�P��$���Q��c�BX�H�у�;���1���U��
�H�J�@�B�E_^[���   ;���1����]� ��������������������������������������������U����   SVWQ�� ����8   ������Y�M���E�P��$���Q��c�BX�H�у�;��X1���U��
�H�J�@�B�E_^[���   ;��21����]� ��������������������������������������������U���  SVWQ�������A   ������Y�M���E�P�� ���Q��c�BX�H�у�;��0���   ���}�E_^[��  ;��0����]� �����������������������������������U���  SVWQ�������A   ������Y�M���E�P�� ���Q��c�BX�H�у�;��(0���   ���}�E_^[��  ;��	0����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BX�H�у�;��/��_^[���   ;��/����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BX�H�у�;��/��_^[���   ;��/����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BX�H�у�;��.��_^[���   ;��.����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BX�H �у�;��.��_^[���   ;��.����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BX�H8�у�;��-��_^[���   ;��-����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�BX�H(�у�;��-��_^[���   ;��-����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�HD�Q,�҃�;��,��_^[���   ;��,����]� ����������������������������������U����   SVW��@����0   �������j j �EP��c�QD��Ѓ�;��!,��_^[���   ;��,����]������������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;��+���E�     _^[���   ;��+����]��������������������������������������U����   SVW��@����0   �������j j �EP��c�QD��Ѓ�;��1+��_^[���   ;��!+����]������������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;���*���E�     _^[���   ;��*����]��������������������������������������U����   SVW��@����0   �������EPj �MQ��c�BD��у�;��?*��_^[���   ;��/*����]����������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;���)���E�     _^[���   ;��)����]��������������������������������������U����   SVW��@����0   �������j j �EP��c�QD��Ѓ�;��Q)��_^[���   ;��A)����]������������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;���(���E�     _^[���   ;���(����]��������������������������������������U����   SVW��@����0   �������EPj h'  ��c�QD��Ѓ�;��^(��_^[���   ;��N(����]���������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;���'���E�     _^[���   ;���'����]��������������������������������������U����   SVW��@����0   �������j j h�  ��c�HD��҃�;��q'��_^[���   ;��a'����]������������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;��'���E�     _^[���   ;���&����]��������������������������������������U����   SVW��@����0   �������j j h:  ��c�HD��҃�;��&��_^[���   ;��q&����]������������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;��&���E�     _^[���   ;���%����]��������������������������������������U����   SVWQ��$����7   ������Y�M��E�    �E�    �E�Pj�M�� ����u3���E�R��P��q����XZ_^[���   ;��e%����]Ð   �q����   �qrp �����������������������������������������U����   SVW��@����0   �������j j h�F ��c�HD��҃�;���$��_^[���   ;���$����]������������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;��r$���E�     _^[���   ;��Y$����]��������������������������������������U����   SVW��@����0   �������j j h�_ ��c�HD��҃�;���#��_^[���   ;���#����]������������������������������U����   SVW��@����0   �������E�Q��c�B@�HH�у�;��#���E�     _^[���   ;��i#����]��������������������������������������U����   SVWQ��$����7   ������Y�M��} u3��(�E�    �E�E�E�Pj�M�������u3���   R��P�\t�M��XZ_^[���   ;���"����]�    dt����   ptrp ���������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�QD�BL�Ѓ�;��?"��_^[���   ;��/"����]����������������������������U����   SVW��@����0   ������E�M��E�M�H�EPj�MQ�)����_^[���   ;��!����]����������������������������U����   SVW��@����0   ������   _^[��]�����������������������U����   SVW��(����6   ������} t�E�8 t�E� �Pj�EP�CA�����E��}� u3��5�M������E�}� u3�� �} t�E�M��E�M;H~3���E�_^[���   ;��� ����]������������������������������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;��a ��_^[���   ;��Q ����]������������������������������U����   SVW��@����0   �������EP��c�Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��(����6   ������} u3��m�EP�#�����E��}� u3��T��E��M��I �PP��;��h���E�}� uh0W��C��P�����3����E�M�I ���   ��;��+��_^[���   ;������]��������������������������������������������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M��E����M��B��;��g��_^[���   ;��W����]��������������������U����   SVWQ��4����3   ������Y�M��E����M��B��;����_^[���   ;�������]��������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M��E����M��B��;��g���M��A�E����M��   _^[���   ;��A����]� ���������������������������U����   SVWQ��4����3   ������Y�M��E����M��B��;������M��A�E����M��   _^[���   ;�������]� ���������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ������9   ������Y�M��E�E�}� t�E��U�<� u3��W�E����M��B��;��I��P�M�3���E���j �E��U��P�M�Q�U���M��P��;������u3���   _^[���   ;�������]� ��������������������������������������������������U����   SVWQ������:   ������Y�M��E�E�}� t�E��U�<� u3��G�E��U��P�M����M��B��;��]��P������;+��P�M����������'���   _^[���   ;��(����]� ��������������������������������������������������U����   SVWQ������9   ������Y�M��E��x�u3��   �E��x t�E��@�   �E�    h�F �*7�����E���E�P�P
�����E��}� t8�M��A���E�E����M��B��;��Z���M�9u�E��M�H�E��$�h0W��C��P�������E��@����3�_^[���   ;������]��������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�h0W��C��P�i����3�_^[���   ;������]� �������������������������������U����   SVWQ��$����7   ������Y�M��E����M��B��;��'��9Eu�} u�   �<�EP�MQ��(�����(��P�M�����(����J%���M�*����t3���   _^[���   ;�������]� ���������������������������������������������������U����   SVWQ��4����3   ������Y�M��E� �������_^[��]� ����������������������U����   SVWQ��4����3   ������Y�M��E� �������_^[��]� ����������������������U����   SVWQ��4����3   ������Y�M��E� �������_^[��]� ����������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U���  SVW��������   ������} u3��  �E���M�B��;�����E�j h@  ������P�2�����E�������E������ǅ�������E������ǅ����:�ǅ����۽ǅ����܊ǅ ����ǅ�����ǅ�����ǅ�����ǅ����ǅ����ǅ����ǅ �����ǅ$���-�ǅ(���+�ǅ,����ǅ0����ǅ4���(�ǅ8�����ǅ<����ǅ@����ǅD�����ǅH�����ǅL�����ǅP���l�ǅT���!�ǅX����ǅ\���q�ǅ`���    ǅd���    ǅh���׊ǅl���&�h@  ������P�MQ�U�Rj�"4����R��P�0��y��XZ_^[��  ;�������]Ë�   8�����@  D�np �����������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��W,���E�� �W�E��M�H�E��M�H�E�_^[���   ;�������]� ���������������������������������U����   SVWQ��4����3   ������Y�M��M��;����E��t�E�P�-�����E�_^[���   ;��~����]� ������������������������U����   SVWQ��4����3   ������Y�M��M���2��_^[���   ;��%����]������������������U����   SVWQ��4����3   ������Y�M��E��P�E��H��I �Rd��;�����_^[���   ;�������]�����������������������������U����   SVWQ��4����3   ������Y�M��E��P�E��H��I �R\��;��`��_^[���   ;��P����]�����������������������������U����   SVWQ��4����3   ������Y�M���EP�M��Q�E��H�I �Rh��;�����_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U��B�M��Q�J ���   ��;�����_^[���   ;�������]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��B�M��Q�J ���   ��;��e��_^[���   ;��U����]� �������������������������������U���  SVW��l����e   ������} u3��   �E���M�B��;������E�j h�   ��0���P������E��P����E��0���ǅ4������E��p���ǅt���۽ǅx���܊ǅ|���:��E����E���E���h�   ��0���P�MQ�U�Rj�k.����R��P������XZ_^[�Ĕ  ;��?����]ÍI    ��0����   ��np ��������������������������������������������������������������������������������̋�`<����������̋�`L����������̋�`\����������̋�`l����������̋�`����������̋�` ����������̋�`0����������̋�`@����������̋�`P����������̋�`p����������̋�`����������̋�`$����������̋�`4����������̋�`D����������̋�`T����������̋�`d����������̋�`t����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`H����������̋�`X����������̋�`h����������̋�`x����������̋�`����������̋�`����������̋�`,�����������U���,  SVWQ�������K   ������Y�M��}}�B  �E�E��E������E�E���EE�EȋE����EE�E��}�~�E���E�E�+E�E��1�EP�M�Q�U�R�M�����E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;���
����}�Eԃ��EԋE��E���E�P�M�Q�U���M����;���
����}�EP�M�Q�U�R�M��������U��������_^[��,  ;��
����]� ����������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et.�E���E�M��U�E���E�M�U���E�M���_^[��]� ��������������������������������U���8  SVWQ�������N   ������Y�M��E���Eȃ}}�B  �E�E��E������E�E���EE�E��E����EE�E��}�~�E���E�E�+E�E��1�E�P�M�Q�U�R�M��-����E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;��^����}�Eԃ��EԋE��E���E�P�M�Q�U���M����;��.����}�E�P�M�Q�U�R�M��X������U��������_^[��8  ;�������]� ������������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et4�E���E�Mf�f�U�E���E�M�Uf�f��Ef�M�f���_^[��]� ������������������������������������������U���8  SVWQ�������N   ������Y�M��E���Eȃ}}�B  �E�E��E������E�E���EE�E��E����EE�E��}�~�E���E�E�+E�E��1�E�P�M�Q�U�R�M������E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;������}�Eԃ��EԋE��E���E�P�M�Q�U���M����;��}����}�E�P�M�Q�U�R�M���������U��������_^[��8  ;��G����]� �����������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et.�E���E�M��U�E���E�M�U���E�M���_^[��]� ��������������������������������U����   SVWQ��4����3   ������Y�M��E��u�EP�MQ�UR�M��#���83��} ����t�EP�MQ�UR�M��
�����EP�MQ�UR�M����_^[���   ;������]� �������������������������������������������������U���  SVWQ�������E   ������Y�M��} t�} t�} t�} u3��  �Ek� E�E���E�P�MQ�U���M����;�����Eȃ}� u
�E���   ��}� }3���   �E�   �E���E��E�;E���   �E�E����EԋE�E�E�E���E�P�MQ�U���M����;�����Eȃ}� uP�}� ~C�Eԃ��EԋE�E�E�E���E�P�MQ�U���M����;��R����t�
��E��E�뷋E��#��}� }�Eԃ��E��	�Eԃ��E��G���3�_^[��  ;��
����]� ����������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��M����_^[���   ;��� ����]������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E�M�P;QuKjj�M��w����u�   �E���U���E���U�B�A�E���U�B�A�E��H�   �Tjj�M��,����u�B�E���U���E���U�B�A�E���U�B�A�E���U�B�A�E��H�   �E�_^[���   ;��������]� ��������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �EP�M������E�_^[���   ;�������]� ���������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��{���E�_^[���   ;�������]� ������������������������U����   SVWQ������<   ������Y�M��M�����} ��   h�W��C��Phi3ɋE�   �������Q�|$����������E��������E��8 u3��   �} tyh�W��C��
Phi3ɋE�   �������Q�'$������ ����E��� ����H�E��x u/�E��8 t�E����,�����,���R������E��     3���E��M�H�E��M�H�   �3�_^[���   ;��b�����]� ��������������������������������������������������������������������������������������������U����   SVWQ������9   ������Y�M��E��8 t�E���� ����� ���R�������E��     �E��x t�E��H��,�����,���R������E��@    �E��@    �E��@    _^[���   ;��`�����]���������������������������������������������U����   SVWQ������9   ������Y�M��M�����} �5  �E�8 �)  �E�x �  h�W��C��Phi3ɋU�B�   �������Q� "������ ����E��� �����E��8 u3���   �E�x tb�E�x tYh�W��C��
Phi3ɋU�B�   �������Q�!������,����E���,����H�E��x u�M�����3��d�E��M�Q�P�E��M�Q�P�E��H��Q�U��P�M�R�|������E��x t �E��H��Q�U��BP�M�QR�S������   _^[���   ;�������]� �����������������������������������������������������������������������������������������������������������U����   SVWQ������<   ������Y�M��M�����} ��  �} �w  h�W��C��Phi3ɋE�   �������Q�" ����������E��������E��8 u3��-  �} tj�} tdh�W��C��
Phi3ɋE�   �������Q�������� ����E��� ����H�E��x u�M�����3���   �E��M�H�c�E��@   h�W��C��Phi3ɋU��B�   �������Q�V������,����E���,����H�E��x u�M����3��Z�E��M�H�E��H��Q�U��P�MQ�G������} t�E��H��Q�U��BP�MQ�$�������E��H�U��   _^[���   ;��u�����]� �������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    _^[��]��������������������������������U����  SVWQ�������   ������Y�M����]��E�    j �M��q���j �M��g���j �M��]����E��H�U�<�}���  �} �&  �M������j ��p����(����E���k�U��E��J�MċR�UȍE�P�M���Bk�EP��$���Q���������p����H��t����P��x����E�   �	�E����E��E��H�U�;}y�E�P�M���E���k�MQ��8���R�b������M��P�U��@�E��E�P��p���Q��L���R�l�����P�M������E���p����M���t����U���x����q���Q���$��`��������E��`������d����P��h����H�E�P��t���Q�|�����U��$��
�H�J�@�B�E���.����z�E���ٝ����	�E�ٝ����E���.����z�E���ٝ����	�E�ٝ���م���م�����������   �E���.����z�E���ٝ����	�E�ٝ����E���.����z�E���ٝ����	�E�ٝ���م���م�����������   �E��$PQ���$Q���$Q���$����������P������Q��������U����
�H�J�@�B�E��P�M��$Q������R�������M�����P�Q�@�A�]  �E���.����z�E���ٝ����	�E�ٝ����E���.����z�E���ٝ����	�E�ٝ���م���م���������zQ���$Q���$Q���$���������P�E��$P������Q�������U����
�H�J�@�B�E��P�M��$Q������R��������M�����P�Q�@�A�}Q���$Q���$Q���$�� ������P�E��$P�����Q�������U����
�H�J�@�B�E��$P�M��Q��(���R�Y������M�����P�Q�@�A�EP��<���Q��������   ���}��E�    �	�E����E��E�;E}�E��H�U��E���E��ۋE���Uԋ�k�EP�MQ��t���R�8������M��P�Uċ@�EȋE���UԋD�k�EP�MQ������R�������M��P�U��@�E��E�    �	�E����E��E��H�U�E�;���   �E����M��I�u��<�UԋE����k�UR�EP������Q�������U��H�M��P�U��E�P�M�Q�U�R�	  ���E��]�E��E��M��MċU��UȋE��E��M��M��U��U��V����E�R��P��������XZ_^[���  ;��{�����]� �   ������   ������   ������   ������   ��p���   �prev n v3 v2 v1 ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVW��4����3   ������E� �M�I�U�B�E���ٝ<���م<���Q�$�M�A�U�
�E� �M�I��ٝ8���م8���Q�$�U�B�E�H�M�A�U�J��ٝ4���م4���Q�$�M�����E_^[���   ;�������]����������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E�� �M��U���E��@�M�A�U��Z�E��@�M�A�U��Z�E�_^[��]� ������������������������������U����   SVW��4����3   ������E�@�M�aٝ<���م<���Q�$�U�B�E�`ٝ8���م8���Q�$�M��U�"ٝ4���م4���Q�$�M�~���E_^[���   ;��E�����]��������������������������������������������������U���  SVW�������A   ������j �M�����E�@�M�I,�U�B(�E�H ��M�I�U�B(�E�H�M�A�U�J,��E�H���M�A�U�J �E�@�M�I��U�J$���]��E���.����Dz�M�����E�u  �E������]��E�@�M�I,�U�B(�E�H��M�I�U�B�E�H�M�A�U�J ��E�H$���M�A(�U�J �E�@�M�I,��U�
���M��]̋E�@�M�I�U�B�E�H��M�I$�U�B�E�H,�M�A(�U�J��E����M�A(�U�J�E�@�M�I,��U�J���M��]ЋE�@�M�I�U�B�E�H ��M�	�U�B �E�H�M�A�U�J��E�H���M�A�U�J�E�@�M�I��U�J���M��]ԋE�@�M�I,�U�B(�E�H ���M��]؋E�@(�M�I�U�B�E�H,���M��]܋E�@�M�I �U�B�E�H���M��]��E�@ �M�I$�U�B,�E�H���M��]�E�@,�M�I�U�B�E�H$���M��]�E�@�M�I�U�B �E�H���M��]�E�@�M�I(�U�B$�E�H���M��]��E�@$�M�I�U�B�E�H(���M��]�E�@�M�I�U�B�E�H���M��]��   �ű}�ER��P�\��N���XZ_^[��  ;��������]ÍI    d�����0   p�mi �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M�������EP�M��������EP�M��������EP�M���$�����E�_^[���   ;��a�����]� �������������������������������������������U����   SVW��<����1   ������E�@�M�a�U�
�E�@�M�a�U�
���E�@�M�a�U�
��ٝ<���م<���_^[��]�����������������������������������������U����   SVW��4����3   ������j�K   ���E��}� u3���E���H��;��Z���_^[���   ;��J�����]�����������������������U����   SVW��@����0   ������hxh�EPh_� ������_^[���   ;��������]�������������������������U����   SVW��(����6   ������E�8 u�>j�q������E��}� u�)�E��M��E�P�M��Q�҃�;��s����E�     R��P�ܰ�����XZ_^[���   ;��I�����]Ð   �����   �i ����������������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3����EP�U�M��B��;�����_^[���   ;�������]� �������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3����EP�U�M��B��;�����_^[���   ;�������]� �������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3�� ��EP�MQ�UR�E�M��P��;��}���_^[���   ;��m�����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�j��������E�}� t	�E�x u3����EP�U�M��B��;������_^[���   ;��������]� �������������������������������U����   SVWQ��(����6   ������Y�M�j �V������E�}� t	�E�x  u3����EP�U�M��B ��;��U���_^[���   ;��E�����]� �������������������������������U����   SVWQ��(����6   ������Y�M�j$��������E�}� t	�E�x$ u2����EP�U�M��B$��;������_^[���   ;�������]� �������������������������������U����   SVWQ��(����6   ������Y�M�j(�6������E�}� t	�E�x( u3����E�M��P(��;��9���_^[���   ;��)�����]��������������������������������������U����   SVWQ��(����6   ������Y�M�j,�������E�}� t	�E�x, u3����E�M��P,��;�����_^[���   ;�������]��������������������������������������U����   SVWQ��(����6   ������Y�M�j0�������E�}� t	�E�x0 u3����EP�U�M��B0��;�����_^[���   ;�������]� �������������������������������U����   SVWQ��(����6   ������Y�M�j4�������E�}� t	�E�x4 u������EP�MQ�U�M��B4��;�����_^[���   ;��p�����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�j8��������E�}� t	�E�x8 u3����E�M��P8��;������_^[���   ;��������]��������������������������������������U����   SVWQ��(����6   ������Y�M�j<�V������E�}� t	�E�x< u���EP�U�M��B<��;��W���_^[���   ;��G�����]� ���������������������������������U����   SVWQ��(����6   ������Y�M�j@��������E�}� t	�E�x@ u���EP�U�M��B@��;������_^[���   ;�������]� ���������������������������������U����   SVWQ��(����6   ������Y�M�jD�6������E�}� t	�E�xD u3����EP�U�M��BD��;��5���_^[���   ;��%�����]� �������������������������������U����   SVWQ��(����6   ������Y�M�jH�������E�}� t	�E�xH u���EP�U�M��BH��;�����_^[���   ;�������]� ���������������������������������U����   SVWQ��(����6   ������Y�M�jL�������E�}� t	�E�xL u3����E�M��PL��;�����_^[���   ;��	�����]��������������������������������������U����   SVWQ��(����6   ������Y�M�jP�������E�}� t	�E�xP u���E�M��PP��;�����_^[���   ;��{�����]����������������������������������������U����   SVWQ��(����6   ������Y�M�jT��������E�}� t	�E�xT u���E�M��PT��;������_^[���   ;��������]����������������������������������������U����   SVWQ��(����6   ������Y�M�jX�f������E�}� t	�E�xX u���E�M��PX��;��k���_^[���   ;��[�����]����������������������������������������U����   SVWQ��(����6   ������Y�M�j\��������E�}� t	�E�x\ u3����EP�MQ�U�M��B\��;������_^[���   ;��������]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j`�6������E�}� t	�E�x` u3����EP�MQ�U�M��B`��;��1���_^[���   ;��!�����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jd�������E�}� t	�E�xd u�(��EP�MQ�UR�EP�MQ�U�M��Bd��;�����_^[���   ;��w�����]� ���������������������������������U����   SVWQ��(����6   ������Y�M�jh��������E�}� t	�E�xh u3�� ��EP�MQ�UR�E�M��Ph��;������_^[���   ;��������]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�jl�V������E�}� t	�E�xl u3����EP�MQ�U�M��Bl��;��Q���_^[���   ;��A�����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jp�������E�}� t	�E�xp u3����EP�MQ�U�M��Bp��;�����_^[���   ;�������]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jt�������E�}� t	�E�xt u3����EP�MQ�U�M��Bt��;�����_^[���   ;�������]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jx�v������E�}� t	�E�xx u3����EP�U�M��Bx��;��u���_^[���   ;��e�����]� �������������������������������U����   SVWQ��(����6   ������Y�M�j|��������E�}� t	�E�x| u3����EP�MQ�U�M��B|��;������_^[���   ;��������]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �C������E�}� t�E샸�    u����/��EP�MQ�UR�EP�MQ�UR�E�M����   ��;��'���_^[���   ;�������]� �������������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u����/��EP�MQ�UR�EP�MQ�UR�E�M����   ��;��g���_^[���   ;��W�����]� �������������������������������������������������U���p  SVWQ�������\   ������Y�M��M�������E�    �	�E؃��E؋E��M�;H�  �E���U؍�������u�ҋE���U؍�������E�E̋E̋M̋P;Qul�E̋k�MQ�ŰBk�EP������Q�q�����P�Űk�EP�M̋Qk�UR������P�H�����P������Q�m�����P�M������k�E̋k�MQ�ŰBk�EP������Q������P�ŰBk�EP�M̋Qk�UR������P�������P������Q� �����P�M�读��������E�P�MQ�\������ER��P����
���XZ_^[��p  ;�������]� �   ������   ��v ��������������������������������������������������������������������������������������������������������������������������U���  SVWQ�������B   ������Y�M��M������E�    �	�Eȃ��EȋE��M�;H��   �E���Uȍ��������u�ҋE���Uȍ��������E�E��E��k�MQ�M��Y����E��Hk�MQ�M��D����E��Hk�MQ�M��/����E��M��P;Qt�E��Hk�MQ�M������S����EP�MQ�M��;���R��P�H��a���XZ_^[��  ;��������]�    P�����   \�mm ���������������������������������������������������������������������������������U����   SVWQ������=   ������Y�M��M��/����M����$���Q�xM�$����������E�������������P������HQ�tM�$��$��������E�����$������(����P��,����H�E��@    �E�_^[���   ;�������]���������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x ��   �E� �M��������Au
�E��M���E�@�M��A������Au�E��M�A�X�E�@�M��A������Au�E��M�A�X�E� �M��A������z�E��M��X�E�@�M��A������z�E��M�A�X�E�@�M��A������z�E��M�A�X�<�E�M������P�Q�@�A�M����U����A�B�I�J�E��@   _^[��]� �����������������������������������������������������������������������������������������U���  SVWQ�������G   ������Y�M��E��x tvQ�X�$�E���P�M�Q�����R�������P��$���P�������M���P�Q�@�A�EP�M���Q������R�e������M���P�Q�@�A�DQ���$������������E��������� ����P������H�U�E�
��J�H�R�P_^[��  ;��������]� ��������������������������������������������������������������������U����   SVW��4����3   ������E�@�Mٝ<���م<���Q�$�M�A�Mٝ8���م8���Q�$�U��Mٝ4���م4���Q�$�M�f����E_^[���   ;��-�����]������������������������������������������U����   SVW��4����3   ������E�@�M�Aٝ<���م<���Q�$�U�B�E�@ٝ8���م8���Q�$�M��U�ٝ4���م4���Q�$�M�����E_^[���   ;��u�����]��������������������������������������������������U����   SVWQ������9   ������Y�M��E�    �E��x|�E��8 u3��?�E�    �	�E����E��E��M�;H}�E���U����������t	�E���E��͋E�_^[���   ;�������]�����������������������������������������������U����   SVWQ��4����3   ������Y�M��E�� %    _^[��]�����������������������������U����   SVWQ��(����6   ������Y�M��E�E��	�E���E�E��M�;H}!�E���U���������t�E�+E����˃��_^[���   ;�������]� ���������������������������������������U����   SVWQ��(����6   ������Y�M��} |�E��8 u����<�E�    �	�E���E�E��M�;H}�E���U������;Eu�E���Ѓ��_^[���   ;�������]� ����������������������������������������U����   SVWQ������9   ������Y�M��E� �E�    �	�E����E��E��M�;H}0�E���U��������;Eu�]�E���U���蹴��؈]���E���_^[���   ;��V�����]� ������������������������������������������������U����   SVWQ��(����6   ������Y�M��M������E�}��u3��
�   �M���_^[���   ;��������]���������������������������U����   SVWQ��4����3   ������Y�M��E����   @t�����E�� %���3ҹ   ���_^[��]��������������������������������U����   SVWQ������9   ������Y�M��E�    �E�    �	�E����E��E��M�;H} �E���U����������t	�E���E��̋E�_^[���   ;��������]�����������������������������������U����   SVWQ������9   ������Y�M��E�    �E�    �	�E����E��E��M�;H}�E���U���������t	�E���E��͋E�_^[���   ;��'�����]������������������������������������U����   SVWQ������<   ������Y�M��E�    �	�E���E�E��M�;H}�E���U��%����M���M�����E�    �	�E���E�E��M�;H}{�E���U��%   �ud�E���U��������EԋE���E��	�E����E��E��M�;H}2�E���U�������;E�u�E���U���   ��M���M�����q���_^[���   ;��������]������������������������������������������������������������������������U����   SVWQ��$����7   ������Y�M��M��������E�E�M�������$�����$�������$�����$���w}��$����$�`��E� ����E� ����\�E�M���E�M�Q��E�E�M�Q��E�M�Q��-�E�M�Q��E�M�Q���E�M�Q��E�M��_^[���   ;��������]� �I ������2�����������������������������������������������������������������������������U����   SVWQ������9   ������Y�M��M�袿���E�M��Ŀ���E��E;E�t	�}���u�E;E�t	�}���u�^�}���t�E�E��}���t�E�E�}��t�E�M����E����   �ыE����E���   @�M����   �M��_^[���   ;�������]� ���������������������������������������������������������������U����   SVW��@����0   �����󫡨c�H\����;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������E�Q��c�B\�H�у�;������E�     _^[���   ;�������]��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q\�B�Ѓ�;��/���_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q\�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q\�B�Ѓ�;��O���_^[���   ;��?�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B\�H�у�;��ۿ��_^[���   ;��˿����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H\�Q�҃�;��X���_^[���   ;��H�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B\�H�у�;��۾��_^[���   ;��˾����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q\�B �Ѓ�;��_���_^[���   ;��O�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B\�H$�у�;�����_^[���   ;��۽����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H\�Q(�҃�;��h���_^[���   ;��X�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q\�B,�Ѓ�;�����_^[���   ;��Ӽ����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B\�H4�у�;��k���_^[���   ;��[�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B\�HD�у�;�����_^[���   ;��ۻ����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B\�HH�у�;��k���_^[���   ;��[�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q\�B8�Ѓ�;�����_^[���   ;��ߺ����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H\�Q<�҃�;��x���_^[���   ;��h�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B\�H@�у�;������_^[���   ;�������]� �������������������������������������U����   SVWQ������?   ������Y�M�j �M贶���M��}����EȋE�P�M蝶���E�    �	�E���E�E�;E�}.�E�P�M�Q�U�R�M��[����E�P�M�c����E�P�M�W�����R��P��薬��XZ_^[���   ;�������]� �   �����   6�����   4�b a ��������������������������������������������������������U���  SVWQ�������B   ������Y�M��E�P�M莦���}� |o�M��\����E�P�M�t����}� tU�E�    �	�E����E��E�;E�};�E�P�M�H����E�P�M�<����	�Eȃ��EȋE�;E��E�P�M��K�����봸   R��P�@��i���XZ_^[��  ;�������]�    H�����   ������   |�����   z�����   x�b a cnt level ��������������������������������������������������������������������������U����   SVW��@����0   �����󫡨c�H����;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������E�Q��c�B�H�у�;�貶���E�     _^[���   ;�虶����]��������������������������������������U����   SVW��@����0   �������E�Q��c�B�H�у�;��2����E�     _^[���   ;�������]��������������������������������������U����   SVWQ������:   ������Y�M���h�  �E�P��(���Q��c�B���   �у�;�蠵���������������(�������������_^[���   ;��r�����]�����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q�B�Ѓ�;������_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B���   �у�;�舴��_^[���   ;��x�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R��c�H���   �҃�;������_^[���   ;�������]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��c�B�Hx�у�;��o���_^[���   ;��_�����]� �������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q�B$�Ѓ�;������_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q�B�Ѓ�;�胲��_^[���   ;��s�����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q�B �Ѓ�;�����_^[���   ;�������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��c�B�H(�у�;�����_^[���   ;��o�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H�Q,�҃�;�����_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��c�Q�B0�Ѓ�;�胰��_^[���   ;��s�����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��c�B�H<�у�;������_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P��c�Q���   �Ѓ�(;��h���_^[���   ;��X�����]�$ ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��c�B�H@�у�;��߮��_^[���   ;��Ϯ����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M��̽����P�M��n�����Pj j �E�P��c�Q�BH�Ѓ� ;��G���_^[���   ;��7�����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q�B�Ѓ�;��ϭ��_^[���   ;�迭����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q�B�Ѓ�;��_���_^[���   ;��O�����]����������������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M�Q��c�B�HH�у� ;��Ӭ��_^[���   ;��ì����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H�QX�҃�;��X���_^[���   ;��H�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H\�у�;��۫��_^[���   ;��˫����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q�Bl�Ѓ�;��_���_^[���   ;��O�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q�Bp�Ѓ�;�����_^[���   ;��ߪ����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�Ht�у�;��{���_^[���   ;��k�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H���   �҃�;������_^[���   ;�������]� �������������������������������U����   SVWQ��$����7   ������Y�M���EP�MQ�U�R��(���P��c�Q���   �Ѓ�;��m���P�M�ש����(���赶���E_^[���   ;��F�����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q���   �Ѓ�;��ܨ��_^[���   ;��̨����]�������������������������U����   SVW��@����0   �����󫡨c�H����;��}���_^[���   ;��m�����]��������������������������U����   SVW��@����0   �������E�Q��c�B�H�у�;������E�     _^[���   ;��������]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR�E�P��c�Q�B�Ѓ�;��w���_^[���   ;��g�����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��c�B�H�у�;������_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��c�Q�B�Ѓ�;�����_^[���   ;��o�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��c�H�Q�҃�;�����_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M��n������M��d����H �G@��;��~���_^[���   ;��n�����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M��ޑ�����M��ԑ���H �GD��;�����_^[���   ;��ޤ����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��M��\����xH u3��#�M��J������M��@������H �FH��;��X���_^[���   ;��H�����]�������������������������������������U����   SVWQ��4����3   ������Y�M��M��̐���xL u3��/��EP�MQ�UR�M�謐�����M�袐���H �GL��;�輣��_^[���   ;�謣����]� ��������������������������������������U���  SVWQ�������D   ������Y�XD3ŉE��M�} t<�M�������E�P�M��������M������H �WL��;������M��M��g����} t?�������>���P�M�6����������[����M�軏���@@�Ẽ}� t�E�P�M����R��P����.���XZ_^[�M�3�������  ;�衢����]� �I    ������   ��bc �����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��������M��܎���H �WH��;������_^[���   ;�������]� ��������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��Z������M��P����H �WD��;��j���_^[���   ;��Z�����]� ������������������������������������U����   SVWQ��4����3   ������Y�M��M��܍���xP u������;��EP�MQ�UR�EP�MQ�UR�M�譍�����M�裍���H �GP��;�轠��_^[���   ;�譠����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��M��,����xT u������+��EP�MQ�M��������M������H �WT��;�����_^[���   ;�������]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��M�茌���xX u�'��EP�M��v������M��l����H �WX��;�膟��_^[���   ;��v�����]� ��������������������������������U����   SVW��$����7   ������M��W����E�P�MQ�ϰ������t�}� u3���E�P�M�Q�U�R�E�P�M��R���R��P�T��V���XZ_^[���   ;��Ӟ����]ÍI    \�����   h�dat ����������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �M��A    �U��B    �E��@    �E�_^[��]�����������������������������������U����   SVW��<����1   ������E��<�����<���t��E��h�E��h�   _^[��]� ��������������������������������U����   SVW������:   ������E�����������������������q  ������$�\��   �]  ��h����h�=�h��   �EP耞����=H&  }
������&  �} u
������  hX��C��Phij�������� ����� ��� t�� ����I���������
ǅ���    ������|h�=|h t�EP�|h�$����   �   �EP�MQ�H�������u����   �   �|�U����u��h����hu\�
���蕖���=|h t?�|h��8�����8�����,�����,��� tj��,����+���������
ǅ���    �|h    �   ����_^[���   ;��ɛ����]Ð��������D�������������������������������������������������������������������������������������������������������������������������������U����   SVW��4����3   ������j�   ���E��}� t	�E��x u����0��E P�MQ�UR�EP�MQ�UR�EP�M��Q�҃�;������_^[���   ;�豚����]����������������������������������������������U����   SVW��@����0   ������h�h�EPh�f �԰����_^[���   ;��<�����]�������������������������U����   SVW������?   ������j�{������E��}� t	�E��x uǅ��������M�q���������E�E8P�M4Q�U0R�E,P�M(Q���̍UR�8����EP�M��Q�҃�4������M�*��������R��P�������XZ_^[���   ;��f�����]Ë�   ������   ��_$ArrayPad �����������������������������������������������������������������U����   SVW��4����3   ������j�[������E��}� t	�E��x u3����EP�MQ�U��B�Ѓ�;�覘��_^[���   ;�薘����]�����������������������������������U����   SVW��4����3   ������j��������E��}� t	�E��x u3����EP�M��Q�҃�;�����_^[���   ;��
�����]��������������������������������������̋�U����M�h�C�X���u/�E�    �	�E����E��}�}�M�k����hQ�w������ڋE���]��������������������������������̋�U����M�h�C�\���}/�E�    �	�E����E��}�}�M�k����hQ�θ�����ڋ�]�������������������̋�U��Qh�C�X���u/�E�    �	�E����E��}�}�M�k����hQ謢�����ڋ�]������������������������̋�U��Qh�C�\���}/�E�    �	�E����E��}�}�M�k����hQ�������ڋ�]������������������������̋�U��Q�M��E��     h�h�,������E���]����������̋�U��Q�M��E��M��U��:}�E��k����hQ�������E���]� ����������������������̋�U��Q�M��E��8}�M��k��hR�G�������]��������������������̋�U��h�h�y�����]������������̋�U��E���M��U�k��hP�E�����]������������������������̋�U��E�k����hQ賲����]������������������̋�U��E��k��hP�ߡ����]������������������̋�U��E��k��hP�S�����]������������������̋�U��Qj 芢����芽����@P�EP�=������} t�M�M���E�hX�`�����@P�U�R�������K�����@Ph �������X�����]����������������������������������̋�U��EPj �MQ�URj��������u�]�����������̋�U��EP�MQ�UR�Ϙ����]���������������������̋�U��E��M�B��PhtX�i�����]��������������̋�U����EP�MQ�U�P�MQ������E��}� uJ� i��u$� i��� i�i裂��h0�蕮����hi�M������h<��M�Q�J����E���]������������������������������������̋�U��Q�M�jh�C�M�莟���E�� �"�E���]������������������������̋�U��EP�MQ�UR�EP�j�����]�����������������̋�U��E�Q�UR�Ց����]�������̋�U��EP�MQ�UR�EP�	�����]�����������������̋�U�츄X]����̋�U��j�h��d�    P��L�XD3�P�E�d�    h�X�M��&����E�    �E�P�M��G���h���M�Q������E������M�螐���M�d�    Y��]�����������������������������̋�U��j�h�d�    P��L�XD3�P�E�d�    h�X�M�薜���E�    �E�P�M��E���h@"�M�Q�j����E������M������M�d�    Y��]�����������������������������̋�U��Q�M��EP�M�藧���M���X�E���]� ��������̋�U��Q�M��E�� �X�M�������]������������������̋�U��Q�M��M��w����E��t�M�Q�������E���]� �����������������̋�U��Q�M��EP�M��g����M���X�E���]� ��������̋�U��j�hH�d�    P��L�XD3�P�E�d�    h Y�M��6����E�    �E�P�M��y��h�"�M�Q�
����E������M�讎���M�d�    Y��]�����������������������������̋�U��Q�M��EP�M��7����M�� Y�E���]� ��������̋�U��Q�M��E��  Y�M�责����]������������������̋�U��Q�M��M��z���E��t�M�Q观�����E���]� �����������������̋�U��Q�M��EP�M������M�� Y�E���]� ��������̋�U��} u�EP�MQh�*訓����]��������������̋�U��Q�E�8u�Fj�MQ�d��E��}� u�U�U�   �#�}�u�E�    ��M�9t
j�`����]����������������������̋�U��EP�h�]���������������̋�U��EP�l�]���������������̋�U��EP�p�]���������������̋�U��EP�t�]����������������u�U��� PRSVW�Ej P�-�����_^[ZX��]�����������̋�U��QSVW3���9>�ى}�~B�F�8ǁ|�����u�Pс<����t�F�L8�UQR�X������E�@��;�E�|�_^[��]���������������������������������̋�U��V���t!��tS�]��tW�̋�����F�V�3_[^]� �������������̋�U��QSVW��3���;�tS9>�}�~L��    �F�8Ǻ����9T�u
�@�9t�N�T�ERP葭��������̋E�@��;�E�|������̋u3��ƅ�tV�@G��u���tJ9u9Vu
9Vu9Vt�MWVQ�`���������̋F9T0�t�MWVQ�D���������̋vO��u�_^[��]� ����������������������������������������������������������̀=$i uj jj j j �$i蜓��P�������������������������������jjj j j �l������������������̋�U��QS�E���E�d�    �d�    �E�]�m��c���[��]� ����������������������������XY�$�����������XY�$�����������XY�$����������̋�U���SVWd�5    �u��E��j �EP�M�Q�UR�}����E�H����U�Jd�=    �]��;d�    _^[��]� ����������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�ё���� �E�_^[�E���]���������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ聑���� �E�_^[�E���]���������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�1����� �E�_^[�E���]��������������������̋�U��E�HQ�U�B(Pj �M�QR�,~����]� �����������������������̋�U����E�    �E��XD�M�3��E��U�U�E�E��M���M�d�    �E�E�d�    �UR�EP�MQ��}���E�E�d�    �E��]����������������������������������̋�U��Q��E�H3M����j �MQ�U�BP�M�QRj �EP�M�QR�EP������� �E��E���]��������������������̋�U���8S�}#  u���M��   ��   �E�    �E� �XD�M�3��E��U�U�E�E�M�M�U �U��E�    �E�    �E�    �e�m�d�    �E؍E�d�    �E�   �E�E̋M�M��E������   �UԍE�P�M�R�Uԃ��E�    �}� td�    ��]؉d�    �	�E�d�    �E�[��]��������������������������������������������������������������������̋�U��QS��E�H3M�W����M�Q��ft�E�@$   �   �v�tj�M�QR�E�HQ�U�BPj �MQ�U�BP�MQ�L����� �U�z$ u�EP�MQ�`���j j j j j �U�Rh#  �{�����E��]�c�k ��   [��]���������������������������������������������������̋�U��Q�} �E�HSV�pW�M�����|8����u�t���E��MN��9L���};H~���u�M���ރ} }̋E�M�UF�1�:;xw;�v�St���M�_��^��[��]��������������������������������̋�U��EV�u�� ������   �N�������   ��^]��������������������̋�U���������   ��t�M9t�@��u��   ]�3�]�������������������̋�U��V訩���u;��   u蘩���N���   ^]�臩�����   �x t�H;�t���x u�^]�Us���V�P^]��������������������������;XDu���"�������������������̋�U��蟪���k����,i�} t�m����]�������������̋�U��]���������̋�U���<Iָ�@Iд�DI���HI���LI��PIָ�TI��XI��\I	��`I��]�������������������������������������̋�U��Q�(i�E��M�(i�E���]������������������̋�U��Q�M��EP�M�Q�~������]� ����������������̋�U��Q�M��E�� �Y�M�Q�Р������]��������������̋�U��Q�M��M��As���E��t�M�Q�v�����E���]� �����������������̋�U��Q�M��EP�M�Q蔣������]� ����������������̋�U��Q�M��E�P��������]�������̋�U��Q�M��E���	P�M��	Q�J������������]� �������������������̋�U��Q�M��E���	P�M��	Q�
���������؋�]� ��������������������̋�U��Q�M��E���	P�M��	Q�ʠ����3҅���]� �����������������̋�U��Q�M��E�����]�������������̋�U��Q�M��E�� �Y�E���]� ��������������������̋�U��Q�M��E���]� �������������̃=Py t-U�������$�,$�Ã=Py t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$������������������������������������������������������̋�U��� VW�   ��Y�}��E�E��M�M��} t�U���t�E� @��M�Q�U�R�E�P�M�Q�|�_^��]� ���������������������̋�U��Q�M��E�� �Y�M��A    �U��B    �E���]�������������������̋�U��Q�M��M��>����E��t�M�Q�7s�����E���]� �����������������̋�U����M��E�� �Y�M�9 tJ�U�P���������E��M�Q� ������U��B�E��x t�M�R�E�P�M��QR�0������
�E��@    �M��A   �E���]� ��������������������������������������������̋�U��Q�M��E�� �Y�M��U��A�M��A    �E���]� ���������������̋�U����M��E�� �Y�M��U�B�A�M��y ta�U�z tL�E�HQ���������E��U�R��������M��A�U��z t�E�HQ�U�R�E��HQ�(������
�U��B    ��E��M�Q�P�E���]� ������������������������������������������������̋�U����M��E�;E��   �M��U�B�A�M��y ta�U�z tL�E�HQ�3��������E��U�R�&������M��A�U��z t�E�HQ�U�R�E��HQ�U������
�U��B    ��E��M�Q�P�E���]� ���������������������������������������������̋�U��Q�M��E�� �Y�M��y t�U��BP�݋������]������������������̋�U��Q�M��E��x t
�M��A���Z��]�����������̋�U��Q�M��EP�M�肃���M��$Z�E���]� ��������̋�U��Q�M��M��.t���E��t�M�Q��o�����E���]� �����������������̋�U��Q�M��EP�M��5����M��$Z�E���]� ��������̋�U��Q�M��E�� $Z�M��U�����]������������������̋�U��Q�M��EP�M�貂���M��4Z�E���]� ��������̋�U��Q�M��M��&y���E��t�M�Q��n�����E���]� �����������������̋�U��Q�M��EP�M��e����M��4Z�E���]� ��������̋�U��Q�M��E�� 4Z�M�腌����]������������������̋�U��Q�M��EP�M��in���M��DZ�E���]� ��������̋�U��Q�M��M�聄���E��t�M�Q�'n�����E���]� �����������������̋�U��Q�M��EP�M��pe���M��DZ�E���]� ��������̋�U��Q�M��E�� DZ�M���w����]������������������̋�U��E�4i]�����������������̋�U��Q�4i�E��M�Q�p~�����E��}� t�UR�EP�MQ�UR�EP�U����&j�r�����MQ�UR�EP�MQ�UR��~������]���������������������������������������̋�U���8  �XD3ŉE�ǅ����    jLj ������P�������������M��� ����U��E�    ǅ���    ������������������������������������f������f������f������f������f������f�������������ǅ ���  �E�������M�������U�B�������ǅ���� �ǅ����   �M����������E�j ����U�R������������� u�}� u
j�p����h ����P����M�3�舍����]���������������������������������������������������������������������������������������̋�U��Q�E�    �4i�E��M�Q�9|�����E��UR�m�����E�E�4i�E���]������������������������������̋�U��Q�E�    �4i�E��M�Q��{�����E��E���]���������������������̋�U��EP�MQ�UR�EP�MQ��|����]�������������̋�U��EP�MQ�UR�EP�MQ�|����]�������������̋�U��j�h0#h"�d�    P���SVW�XD1E�3�P�E�d�    �} t�}t	�E�    ��E�   �EԉE܃}� uh@\j jah�[j�<h������u̃}� u.辆���    j jah�[h�[h@\�|��������b  3҃} �U؃}� uhd[j jbh�[j��g������u̃}� u.�Z����    j jbh�[h�[hd[�{���������  j��h�����E�    �<y�M��	�U�B�E�}� t�M�Q;Uu���}��   �}� th�E�H���U�J�E�H�M��}� uH�U�z t�E�H�U���M�9 t�U��M�Q�P��E�H�<yj�U�R�|t�����43�uh�Zj jh�[j��f������u��E������Q����    ��   �}� tr�U�B���M�A�U�B�E��M�;<ytM�U�z t�E�H�U���M��E�H�J�U��    �E�<y�H�<y�E��M�<y�h�   h�Zjj��_�����E�}� u�E�����裄���    �L�U��    �E�<y�H�=<y t�<y�E��M��A   �E�   �U�E�B�M�<y�E������   �j������ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP��q�����E��E�    �E���]�����������������̋�U��EP�MQ�UR�EP�MQ�UR��r����]���������̋�U��X"  �<c���XD3ŉE��E�    �E�    �} u
�   �  3�f������h  ������Qj �����u8j h<  h�[h|bh bh�ah  ������R�L�����P�ln�����������E��M�Q��������@v`�U�R�ԏ�����M��TA��U�j hE  h�[h|bh�`j�EP�M�������+����  +���P�M�Q��n����P��m�����} t'�UR�n�������@v�EP�]������M�TA��U�蕁��� ������舁���     �}uǅ�����_�
ǅ�����_�M���t�E�������
ǅ�����_�M���t�}uǅ����|_�
ǅ�����_�E���tǅ����t_�
ǅ�����_�} t�U�������
ǅ�����_�} tǅ����`_�
ǅ�����_�} t�E�������
ǅ�����_�} tǅ����L_�
ǅ�����_�}� t�M��������'�} t�U�������
ǅ�����_�������������}� tǅ����PZ�
ǅ�����_�} tǅ����4_�
ǅ�����_������Q������R������P������Q������R������P������Q������R������P������Q������R�E�P�M���ZRhh^h�  h   ������P轇����D�E�}� }*j h`  h�[h|bhH^j"j����Q�y\���� �q����������}� }8j hc  h�[h|bh�]h(]h   ������P�6�����P�Vk����h  h�\������Q覄����������������uj�rm����j�,c��������u�   �3��M�3������]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��} u��EP�MQ�UR�EP�MQ�kr����]���������������������̋�U��} t�E;Et�M;Mt�E��U$R�E P�MQ�UR�EP�r�����E]�������������������������������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP��k�����E��E�    �E���]�����������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+��������������������������������������̋�U��j�EP�k����]�����������̋�U����} u3��k  3��} ���E��}� uh�cj j7hcj�?]������u̃}� u0��{���    j j7hch�bh�c�q�����   �  �} t�U;U��   �EPj �MQ�؆����3҃} �U��}� uh�bj j=hcj�\������u̃}� u-�7{���    j j=hch�bh�b�p�����   �~�M;M҃��U�uh�bj j>hcj�T\������u̃}� u-��z��� "   j j>hch�bh�b�,p�����"   ��   ��MQ�UR�EP�ye����3���]������������������������������������������������������������������������������������������������������������̋�U����} u3��@  3��} ���E��}� uh�cj j6h�cj�O[������u̃}� u0��y���    j j6h�ch�ch�c�'o�����   ��   3҃} �U��}� uh�bj j7h�cj��Z������u̃}� u-�ky���    j j7h�ch�ch�b��n�����   �w�M;M҃��U�uh�bj j8h�cj�Z������u̃}� u-�
y��� "   j j8h�ch�ch�b�`n�����"   ��MQ�UR�EP�2c����3���]���������������������������������������������������������������������������������������̃= y ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uZ�zG ��= y t2���\$�D$%�  =�  u�<$f�$f��f���d$u�wy�������$�T$�D$�   ��ÍT$�b����P��<$f�<$t�s����  ��T$��  ���   �~b����   �  ���   �L$���S  ���x����u���=(i ��g���E�   �@z���=(i ��g���E�   �����ZÍT$�b���D$uA�3���   ���D$u����   �3��3�%�� D$uÍT$��a���D$��%  ����� =  �uT$u���u���t��Q���$�\$��q��W����Y�a���t���g���   �B����D$%�� D$������؋D$%���D$t=�f   �l$���D$�   t�-�L��t��   ����������f�����f�������f�����   ��������������-0M�   ���������ٱ ����u�E�������ٛ���u���������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���@�} t�} v	�E�   ��E�    �ẺEԃ}� uh ej j4h�dj�fV������u̃}� u0��t���    j j4h�dhldh e�>j�����   �G  �U� �}�tI�}���t@�}v:�E��9�Hs��H�M��	�U���UȋE�Ph�   �M��Q������3҃} �UЃ}� uhDdj j8h�dj�U������u̃}� u0�-t���    j j8h�dhldhDd�i�����   �   �M�MċUăz |�Eă8 s��s���    �   �a�M�M��U��z|�E��8�o@�v�s���    �   �3�MQ�U�R�j�����E؃}� u�E�P�MQ�UR�E������E؋E؋�]���������������������������������������������������������������������������������������������������������������������������������̋�U���03��} ���Eԃ}� uhDdj j\h�dj�,T������u̃}� u*�r���    j j\h�dhpehDd�h����3��S�U�UЋEЃx |�MЃ9 s�kr���    3��+�UR�E�P�qi�����E؃}� u�M�Q�ˆ������3���]�������������������������������������������������̋�U����E�P����M��� �>ՋU���ޱ�j h��� RQ�o���E��U�}�|	�}��o@�v�E������E������} t�E�M���U�P�E��U��]�������������������������������������������̋T$�L$��ti3��D$��u��   r�=Py t��Y��W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$��������������������������������������̃= y ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�Ij ��= y t2���\$�D$%�  =�  u�<$f�$f��f���d$u�m�����$�Tk���   ��ÍT$�[��R��<$tmf�<$t�jk��=  �?s-����������������=(i �L`���   � E�~d��w8�D$��%�� D$u'��   ���t�������蟂������ u�|$ u����-0M�   �=(i ��_���   � E�`��Z������������������������������������������������������������������������������������������̃��$�/j���   ��ÍT$��Y��R��<$�D$tQf�<$t�Aj���   �u���=(i �1_���   �0E�cc���  �u,��� u%�|$ u��蒁���"��� u�|$ u�%   �t����-0M�   �=(i ��^���   �0E�_��Z������������������������������������������������������̋�U��Q�|sP�6b�����E��}� t�U�j�|����jj ��L�����r����]�����������������̋�U��Q�E�    �|sP��a�����E��MQ�CS�����|s�E���]��������������������������̋�U��|sP�a����]�����������̋�U��j�hP#h"�d�    P���SVW�XD1E�3�P�E�d�    �}�u�=U���     �)m��� 	   ����  �} |�E;�ws	�E�   ��E�    �M؉M��}� uh�fj j/h�fj�CN������u̃}� u9��T���     �l��� 	   j j/h�fhpfh�f�b��������  �E���M������ x�D
������؉E�uh<fj j0h�fj�M������u̃}� u9�HT���     �4l��� 	   j j0h�fhpfh<f�a��������   �UR��I�����E�    �E���M������ x�D
��t�MQ��~�����E��4��k��� 	   �E�����3�uh�ej j:h�fj�M������u��E������   ��MQ�II����ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������̋�U��QV�EP�:V�������t]�}u� x���   ��u�}u(� x�HD��tj��U������j��U����;�t�UR��U����P�����t	�E�    �	����E��EP�fm�����M���U������ x�D �}� t�M�Q��I��������3�^��]����������������������������������������������������̋�U��j�hp#h"�d�    P�ČSVW�XD1E�3�P�E�d�    �E�    3��} ���E��}� uh�hj jYh@hj��J������u̃}� u9�fQ���     �Ri���    j jYh@hh$hh�h�^��������  j0j �UR�t�����}�u�Q���     �i��� 	   ����a  �} |�E;�wsǅ|���   �
ǅ|���    ��|����M��}� uh�gj j]h@hj�J������u̃}� u9�P���     �h��� 	   j j]h@hh$hh�g��]���������  �E���M������ x�D
������؉E�uh`gj j^h@hj�I������u̃}� u9�P���     �h��� 	   j j^h@hh$hh`g�[]��������H  �UR�E�����E�    �E���M������ x�D
��u9�g��� 	   �E�����3�uh�ej jgh@hj��H������u��  �E���M������ x�
P���%����E܃}��8  �}�t
�}���   �}�u�    �Uf�J��   �Mf�A�U�E��M�U�Q�   �Mf�A3ҋEf�P3ɋUf�J3��Mf�A
�U�B(    �B,    �E�@     �@$    �M�A    �A    �}�u�U�B    �Jj �E�Pj j j �M���U������ x�Q����E��}� t�U�E��B�
�M�A    �  �:�}� u�5f��� 	   �E������q  ����P��E�����E������T  3ҋEf�P3ɋUf�J3��Mf�A
3ҋEf�P�   �Uf�J�E�P�M���U������ x�Q�����u���P�YE�����E�������  �U���t�E�H��$  �Uf�J��E�H�ɶ  �Uf�J�}� u�}� tc�E�P�M�Q�����t�U�R�E�P�����u�E������s  j��M�Q�U�R�E�P�M�Q�U�R�E�P�jZ�����M�A �Q$��U�B     �B$    �}� u�}� tc�E�P�M�Q�����t�U�R�E�P�����u�E�������   j��M�Q�U�R�E�P�M�Q�U�R�E�P��Y�����M�A�Q��U�E�H �J�@$�B�}� u�}� t`�M�Q�U�R�����t�E�P�M�Q�����u	�E������uj��U�R�E�P�M�Q�U�R�E�P�M�Q�lY�����M�A(�Q,��U�E�H �J(�@$�B,�M�UȉQ�E�H�� �  �Uf�J�E�     �M�A    �E������   ��UR�hA����ËE؋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���j �E�P�MQj@�UR�EP�w�����E��}� t	�E�������M��M�E��]�����������������������������̋�U���j �E�P�MQ�UR�EP�MQ�v�����E��}� t	�E�������U��U�E��]���������������������������̋�U���j �E�P�MQj@�UR�EP�w�����E��}� t	�E�������M��M�E��]�����������������������������̋�U���j �E�P�MQ�UR�EP�MQ�v�����E��}� t	�E�������U��U�E��]���������������������������̋�U��Qj �EP�����u����E���E�    �}� t�M�Q��?��������3���]���������������������������̋�U���\  �XD3ŉE�3��} �������������� uh�jj jOh`jj�)A������u̃����� u.�_���    j jOh`jh4jh�j��T��������	  ǅ����   ������ uh�ij jTh`jj��@������u̃����� u.�@_���    j jTh`jh4jh�i�T��������  3��} �������������� uh�ij jUh`jj�T@������u̃����� u.��^���    j jUh`jh4jh�i�)T��������4  ������R�EP����E��}��uq�����������������������������������������w.��������HJ�$�<J�G^���    ��:^���    ��-^���    ����   ��������   ���#������E�������Q�h�����M�A�Q������R�h�����M�A�Q������R�rh�����M�A�Q�U�������B j jwh`jh4jh�h������Qh  �U��$R�_����P�I�����E��M�3��Xb����]ÍI UIbIoI   ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���\  �XD3ŉE�3��}��������������� u!h kj h�   h`jj�=������u̃����� u1�5\���    j h�   h`jh�jh k�Q��������  3҃} ������������ u!h�jj h�   h`jj�C=������u̃����� u1��[���    j h�   h`jh�jh�j�Q��������  ǅ����   ������ u!h�ij h�   h`jj��<������u̃����� u1�T[���    j h�   h`jh�jh�i�P��������1  ������R�EP�����uq�����������������������������������������w.���������M�$��M��Z���    ��Z���    ��Z���    ����   ��������   ���#������E�������Q�%e�����M�A�Q������R�e�����M�A�Q������R��d�����M�A�Q�U�������B j h�   h`jh�jh�h������Qh  �U��$R�[����P�$F����3��M�3���^����]��L�L�L   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�8 u�M�y u�������T�U�R�EP�����t�M�Q�U�R�����u�������(j��E�P�M�Q�U�R�E�P�M�Q�U�R�	N������]����������������������������������������W�|$�n��$    ���L$W��   t�����t=��   u�������~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�����tf�����   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_������������������������������������������������������������������������̋�U����E��}�E��E��}�U��E��U���]����������̋�U���(�E�E��M�M��U�U��}��g  �E��$�DR�M�Q�U�R��  ���E�}� t�E�E��s�M���Q�U���R��  ���E�}� t�E�E��F�M���Q�U���R�  ���E�}� t�E�E���M���Q�U���R�  ���E�E�E�M�M�E���   �U�R�E�P�Y  ���E�}� t�M�M��F�U���R�E���P�2  ���E�}� t�M�M���U���R�E���P�  ���E܋M܉M��E��i�U�R�E�P��   ���E�}� t�M�M���U���R�E���P��   ���E؋E��*�M�Q�U�R�   ���3���EP�M�Q�U�R�  ����]Ð'RR�QjQ�P�����������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U���M��+�P�   ����]�����������������̋�U��} t3��} ���D ��E�E]����������������̋�U����} �R  �EP�MQ�Q	  ���E��}� t�E��O  �U��R�E��P�*	  ���E��}� t�E��(  �M��Q�U��R�	  ���E��}� t�E��  �E��P�M��Q��  ���E��}� t�E���  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q�g  ���E��}� t�E��e  �U��R�E��P�@  ���E��}� t�E��>  �M�� �M�U�� �U�E�� �E�����MM�M�UU�U�E�E��}���  �M��$��Y�U��R�E��P��  ���E��}� t�E���  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q�  ���E��}� t�E��}  �U��R�E��P�X  ���E��}� t�E��V  �M��Q�U��R�1  ���E��}� t�E��/  �E��P�M��Q�
  ���E��}� t�E��  �U��R�E��P��  ���E��}� t�E���  3���  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q�  ���E��}� t�E��  �U��R�E��P�g  ���E��}� t�E��e  �M��Q�U��R�@  ���E��}� t�E��>  �E��P�M��Q�  ���E��}� t�E��  �U��	R�E��	P��  ���E��}� t�E���  �M��Q�U��R��  ���E��}� t�E���  �E��P�M��Q��������  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R�b  ���E��}� t�E��`  �E��P�M��Q�;  ���E��}� t�E��9  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R��  ���E��}� t�E���  �E��
P�M��
Q��  ���E��}� t�E���  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R��  ���  �E��P�M��Q�]  ���E��}� t�E��[  �U��R�E��P�6  ���E��}� t�E��4  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q��  ���E��}� t�E���   �U��R�E��P��  ���E��}� t�E��   �M��Q�U��R�  ���E��}� t�E��   �E��P�M��Q�s  ���E��}� t�E��t�U��R�E��P�o������E��}� t�M��M��F�U��R�E��P�H������E��}� t�M��M���U��R�E��P�!������E��M��M�E��3���]Ë��U�V%XNY�U�V�W*Y�U�V�WYlU�V�W�XEU]V�W�XU6VbW�X�TV;WgX�T�UW@X�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U���M��;�tK�E�E��M�M�U�R�E�P�������E�}� t�M�M���U���R�E��P�\������E�E��3���]�������������������������������������������̋�U��� �E�E��M�M��U��E��
;��   �U�U��E�E�M�Q�U�R��������E�}� t�E�E��s�M���Q�U��R�������E�}� t�E�E��F�M���Q�U��R�������E�}� t�E�E���M���Q�U��R�n������E��E��E�M�M�E��3���]�����������������������������������������������������������������̃= y ��B�����\$�D$%�  =�  u�<$f�$f��f���d$��B��� �~D$f(�kf(�f(�fs�4f~�fT�kf��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�K*�����D$��~D$f��f(�f��=�  |!=2  �fT�k�\�f�L$�D$����f��kfV�kfT�kf�\$�D$�������������������������������������������������������������������������������̃= y ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU险 ��= y t2���\$�D$%�  =�  u�<$f�$f��f���d$u�.�����$�C���   ��ÍT$�2��R��<$tPf�<$t�-��������z�=(i �
8���   �@E�<<���-����������z��������lZ������ u�|$ u����-0M�   �=(i ��7���   �@E�|8��Z���������������������������������������������������������������������������������������̃= y ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�9� ��= y t2���\$�D$%�  =�  u�<$f�$f��f���d$u�M�����$�A���   ��ÍT$�21��R��<$tPf�<$t�-��������z�=(i ��6���   �PE�:���-����������z���������X������ u�|$ u����-0M�   �=(i �56���   �PE��6��Z���������������������������������������������������������������������������������������̋�U��Q�}��   j�!������u3��  �0����u��*��3��  ��5���Ȓ����G���<i��^����}��Y���*��3��U  �2H����|��D����|j �@D������t��V����Y���{*��3��  j�D?�����8i���8i��   �} uW�=8i ~B�8i���8i�=To u��N��j��N������ t�v]���V���RY���	*���3��   �   �}��   �z��h�   h�kjh  j��B�����E��}� tX�U�R�0IP��iQ�!8�����Ѕ�t%j �U�R�?�����Ē�M���U��B�����j�E�P��2����3���3����}u
j �(�����   ��]� ����������������������������������������������������������������������������������������������������������������������̋�U��}u��L���EP�MQ�UR�   ��]� �����������������������̋�U��j�h�#h"�d�    P���SVW�XD1E�3�P�E�d�    �e��E�   �} u�=8i u3��N  �E�    �}t�}uT�=�k t�EP�MQ�UR��k�E�}� t�EP�MQ�UR�DA���E�}� u�E�    �E������E���   �EP�MQ�UR��I���E�}u=�}� u7�EPj �MQ�I���URj �EP��@���=�k t�MQj �UR��k�} t�}u@�EP�MQ�UR�@����u�E�    �}� t�=�k t�EP�MQ�UR��k�E��E������8�E���U��E�P�M�Q�*����Ëe��E�    �E������E��
�E������E�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������̋�U��j�h�#h"�d�    P���SVW�XD1E�3�P�E�d�    �2���E�    �EP�Y   ���E��E������   ��SE��ËE�M�d�    Y_^[��]������������������������������������������̋�U���� yP�44�����E��yQ�"4�����E��U�;U�r�E�+E�����s3��  j�M�Q�O�����E�U�+U���9U���   �}�   s�E�E���E�   �M�M�M�U�;U�r%h�   h lj�E�P�M�Q�8�����E��}� u:�U���U�E�;E�r%h�   h lj�M�Q�U�R�_8�����E��}� u3��W�E�+E����M����U��E��E��M�Q�$����� y�UR�$�����M���U����U��E�P�{$�����y�E��]��������������������������������������������������������������������������������������������������̋�U��EP�T��������؃�]��������������������̋�U��Qh�   h ljjj ��<�����E��E�P�#����� y� y�y�}� u�   ��U��    3���]����������������������̋�U��Qj j j��tP�MQ�.�����E��E���]�������������������������U��WV�u�M�}�����;�v;���  ��   r�=Py tWV����;�^_u^_]������   u������r*��$�tk��Ǻ   ��r����$��j�$��k��$�k��j�j�j#ъ��F�G�F���G������r���$�tk�I #ъ��F���G������r���$�tk�#ъ���������r���$�tk�I kkXkPkHk@k8k0k(k�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�tk���k�k�k�k�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�m�����$��l�I �Ǻ   ��r��+��$�l�$�m�$lHlpl�F#шG��������r�����$�m�I �F#шG�F���G������r�����$�m��F#шG�F�G�F���G�������V�������$�m�I �l�l�l�l�l�l�lm�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�m�� m(m8mLm�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̀�@s�� s����Ë���������������������������̋�U���4�E؉E�3Ƀ} ���Mԃ}� uhmj jph�lj�f������u̃}� u.��8���    j jph�lh�lhm�>.���������   3��} ���EЃ}� uh\lj juh�lj�������u̃}� u.�8���    j juh�lh�lh\l��-��������   �U��B����E��@B   �M��U�Q�E��M��UR�EP�MQ�U�R��P�����E��} u�E��M�E��H���U��J�E��x |!�M��� 3�%�   �E̋M�����E����M�Qj ��-�����E̋E���]����������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR��9����]�������������������̋�U���,�E؉E�3Ƀ} ���Mԃ}� u!hmj h�  h�lj�c������u̃}� u.��6���    j h�  h�lh@mhm�8,��������C�E��@����M��AB   �U��B    �E��     �MQ�UR�EP�M�Q�U���E��E���]����������������������������������������������������̋�U��EPj �MQh[��I����]������������������̋�U��EP�MQ�URh[��jI����]����������������̋�U��EPj �MQh���<I����]������������������̋�U��EP�MQ�URh���
I����]����������������̺`E�,���`E�3���Ƀ=,it����N�������z�����������������̋�U���0  �XD3ŉE��E�    ��E��t
j
�C��������E��}� t
j�r#������E����   ������������������������������������f������f������f������f������f������f�������������ǅ ���  �U�������E�������M�Q�������jPj ������P��?����ǅ����  @�M�������������U� ����E�j ����M�Q���j�V���M�3���8����]�����������������������������������������������������������������������������̋�U��Q��E�E��M��#M��U#Uʉ�E�E���]���������������������̋�U��j�h�#h"�d�    P���SVW�XD1E�3�P�E�d�    3��} ���E؃}� uh\lj j/h�nj�������u̃}� u.�3���    j j/h�nh�nh\l�j(���������  3҃} �Uԃ}� uh�nj j0h�nj�.������u̃}� u.�2���    j j0h�nh�nh�n�(��������  �M�MЋUЋB��@��   �M�Q�rG�����Ẽ}��t!�}��t�U����Ẽ���� x�E���E�PN�MĊQ$������uA�}��t!�}��t�M����Ũ���� x�U���E�PN�E��H$�� ���х�t	�E�    ��E�   �E��Eȃ}� uhpmj j1h�nj�������u̃}� u+�1���    j j1h�nh�nhpm��&���������UR�?�����E�EP��H�����E�    �MQ�p;�����E܋UR�E�Pj�MQ��$�����E��UR�E�P�,�����E������   ��MQ�$����ËE�+E�����M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���E]����̋�U��Q�=�� u���   ��=��}
���   h�   hPojj���P�.�����\y�=\y u?���   h�   hPojj���Q�R.�����\y�=\y u
�   �   �E�    �	�U����U��}�}�E����E�M��\y�����E�    �	�E����E��}�}f�M����U������� x�<�t8�M����U������� x�<�t�M����U������� x�< u�M���ǁ�E�����3���]������������������������������������������������������������������������������������̋�U���)<���Po��t����j�\yQ�a����]�������������������̋�U��}�Er4�}(Hw+�E-�E����P�������M�Q�� �  �E�P��M�� Q�p�]�������������������������������̋�U��}}#�E��P�y�����M�Q�� �  �E�P��M�� Q�p�]�������������������̋�U��}�Er4�}(Hw+�E�H������U�J�E-�E����P�&G������M�� Q�t�]�������������������������������̋�U��}}#�E�H������U�J�E��P��F������M�� Q�t�]�������������������̋�U��j�h�#h"�d�    P���SVW�XD1E�3�P�E�d�    �} uj �  ���@�EP��C�����E�    �MQ�!�����E��E������   ��UR�f����ËE�M�d�    Y_^[��]������������������������������������������̋�U��} uj �n  ���@�EP��'������t����+�M�Q�� @  t�EP��@����P��=��������3�]�����������������������̋�U����E�    �E�E�M�Q����u|�E�H��  tn�U�E�
+H�M��}� ~Z�U�R�E�HQ�U�R�Q@����P�l5����;E�u�E�H��   t�U�B����M�A��U�B�� �M�A�E������U�E�H�
�U��B    �E���]�����������������������������������������������������̋�U��j�   ��]���������������̋�U��j�h$h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    �E�    j�������E�    �E�    �	�E����E��M�;����   �U�\y�<� ��   �M��\y���H��   ��   �U�\y��Q�U�R�9-�����E�   �E��\y���B%�   te�}u%�M��\y��P��������t	�M���M��:�} u4�U�\y���Q��t!�E��\y��R�w�������u�E������E�    �   ��E��\y��R�E�P������������E������   �j��B����Ã}u�E����E܋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������̋�U��Q�EP�MQ�UR��tP�MQ������E��E���]������������������̋�U��j j j�EP�MQ�p����]�������������������̋�U����E�    �E�P�MQ�UR�EP�MQ�UR�D   ���E��}� u�}� t��'����t
��'���M���E���]������������������������̋�U��Q�EP�MQ�UR�EP�MQ�   ���E��}� t�E��3�} u�U�   �E���EP�T@������u�M�   3��룋�]�������������������������̋�U��j j j�EP�[=����]�������̋�U��j�h@$h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    �E�    j�i	�����E�    �=ti vU�ti��9\iu6��+����u!hqj hy  h�pj��������u��\i    ��\i���\i��H�E؃=�H�t�M�;�Hu̃=pI tu�UR�EP�M�Q�UR�EPj j�pI����uP�} t%�MQ�URhTpj j j j ��������u�� h,ph$Uj j j j ��������u��8  �U����  ��t��H��u�E�   �}�v-�MQh pj j j j�������u̋E�    ��  �M����  ��t:�}t4�U����  ��t&�}t h�oh$Uj j j j�:������u̋M��$�MԋU�R�)�����E܃}� u�E�    �r  ��H����H�}� tI�U��    �E��@    �M��A    �U��B�����E܋M�H�U��B   �E��@    �   ���+Ti;Mv�TiU�Ti�
�Ti�����liE�li�li;`iv�li�`i�=di t�di�M܉H�	�U܉Xi�E܋di��U��B    �E܋M�H�U܋E�B�M܋U�Q�E܋M�H�U܋E؉B�M܉dij��HR�E܃�P�&/����j��HQ�U�E܍L Q�	/�����UR��HP�M܃� Q��.�����U܃� �U��E������   �j�<=����ËE��M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�P�MQ�UR�EP�MQ�8������E��}� u�}� t�""����t
�"���U���E���]����������������������������̋�U����} vk�����3��u;E����E�u!hdqj hH  h�pj�������u̃}� u-�!���    j hH  h�ph<qhdq������3��K�U�U�U�EP�MQ�UR�EP��tQ�UR�������E��}� t�EPj �M�Q�,�����E���]��������������������������������������������������������̋�U����E�    �E�P�MQ�UR�EP�MQ�UR�|-�����E��}� u�}� t� ����t
� ���M���E���]������������������������̋�U��Qj j j�EP�MQ�UR��������E��E���]����������������������̋�U��j�h`$h"�d�    P���SVW�XD1E�3�P�E�d�    j������E�    j�EP�MQ�UR�EP�MQ�b   ���E��E������   �j�9����ËE�M�d�    Y_^[��]����������������������������������������������̋�U����E�    �E��M��} u�UR�EP�MQ�U�R�������  �} t�}� u�EP�MQ�&����3��  �=ti vV�ti��9\iu6�A$����u!hqj h�  h�pj�S ������u��\i    ��\i���\i��H�U�=�H�t�E�;�Hu̃=pI ty�MQ�UR�E�P�MQ�U�R�EPj�pI����uR�} t%�MQ�URh$uj j j j �k ������u�� h�th$Uj j j j �I ������u�3��  �}��v`�} t)�UR�EP�M�Qh�tj j j j� ���� ��u���E�Ph pj j j j���������u������    3��3  �}th�U����  ��tZ�E%��  ��tM�} t%�MQ�URhHtj j j j��������u�� h�oh$Uj j j j�p�������u��Qj��HR�E�����P��  ����t1�MQh�sj j j j�/�������u�����    3��t  �EP��)������u!h�sj h  h�pj�B�������u̋U�� �U�E�xu�E�   �}� t8�M�y����u	�U�z t!h�rj h  h�pj���������u��d�M�Q����  ��u�E%��  ��u�E   �M�Ti;Qs1�EPh�rj j j j�C�������u��!���    3��  �} t%�U���$R�E�P��������E��}� u3��_  �#�M���$Q�U�R�"�����E��}� u3��:  3�u���H����H�}� u|�=Ti�s9�U�Ti+B�Ti���+Ti;M�v�TiU��Ti�
�Ti�����E��li+H�li�liU��li�li;`iv�li�`i�U��� �U�E��M�;Hv$�U��E�+BP��HQ�U��E�BP�_&����j��HQ�U�U�R�F&�����}� u�E��M�H�U��E�B�M��U�Q�E��M��H�} u/�} u�U�;U�t!h0rj h�  h�pj���������u̋M�;M�t�}� t�E���   �U��: t�E���U��B�A�8�Xi;M�t!h�qj h�  h�pj��������u̋E��H�Xi�U��z t�E��H�U����7�di;M�t!h�qj h�  h�pj�J�������u̋E���di�=di t�di�E��B�	�M��Xi�U�di��M��A    �U��di�E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�    �E�    �} vk�����3��u;E����E�u!h�uj hA  h�pj��������u̃}� u-����    j hA  h�phhuh�u������3��g�U�U�U��} t�EP������E��MQ�UR�EP�M�Q�UR�L�����E�}� t �E�;E�s�M�+M�Qj �U�U�R�u"�����E��]�����������������������������������������������������������������������̋�U��Qj j j�EP�MQ�1�����E��E���]����������̋�U��j�h�$h"�d�    P���SVW�XD1E�3�P�E�d�    3��} ���E��}� u!h�uj h�  h�pj��������u̃}� u-�!���    j h�  h�ph�uh�u�t����3��c�}�v�����    3��Nj�������E�    j �UR�EP�MQ�UR�EP�7������E��E������   �j�o/����ËE�M�d�    Y_^[��]�������������������������������������������������������������������̋�U��j�EP�T)����]�����������̋�U��j�h�$h"�d�    P��SVW�XD1E�3�P�E�d�    j�������E�    �EP�MQ��(�����E������   �j�.����ËM�d�    Y_^[��]����������������������������������̋�U��Q�=ti vU�ti��9\iu6�����u!hqj h  h�pj��������u��\i    ��\i���\i�} u�l  �}uOj��HP�M�����Q�	  ����t/�URh�zj j j j���������u������    �  �=pI tDj j j �MQj �URj�pI����u%h�zh$Uj j j j ��������u���  �MQ�F ������u!h�sj h%  h�pj��������u̋E�� �E��M��Q����  ��tD�E��xt;�M��Q����  ��t*�E��xt!hHzj h+  h�pj�T�������u̋�H���m  j��HP�M���Q�k  ������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ���oPhxyj j j j�z�����(��u��<�U��� R�E��HQ�U��B%��  ���oQh�xj j j j�<����� ��u�j��HP�M��Q�E��L Q�  ������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ���oPhxj j j j�������(��u��<�U��� R�E��HQ�U��B%��  ���oQhhwj j j j������ ��u̋E��xue�M��y����u	�U��z t!h�vj hd  h�pj��������u̋M��Q��$R��HP�M�Q�n�����U�R�6*�����Q  �E��xu�}u�E   �M��Q;Ut!h�vj hr  h�pj�(�������u̋M��li+Q�li��H����   �M��9 t�U���M��Q�P�6�Xi;E�t!hTvj h�  h�pj���������u̋U��B�Xi�M��y t�U��B�M����5�di;E�t!h vj h�  h�pj�w�������u̋U���di�M��Q��$R��HP�M�Q�B�����U�R�
)�����(�E��@    �M��QR��HP�M��� Q�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�EP�(����]�����������̋�U��j�h�$h"�d�    P���SVW�XD1E�3�P�E�d�    3��} ���E܃}� u!h�uj h�  h�pj�O�������u̃}� u1�����    j h�  h�ph {h�u�$��������8  �=ti vV�ti��9\iu6������u!hqj h�  h�pj���������u��\i    ��\i���\ij��������E�    �UR�������u!h�sj h�  h�pj�w�������u̋M�� �M��U��B%��  ��tC�M��yt:�U��B%��  ��t*�M��yt!hHzj h�  h�pj��������u̋E��xu�}u�E   �M��Q�U��E������   �j�F&����ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������̋�U��Q��H�E��M��H�E���]������������������̋�U��j�h�$h"�d�    P���SVW�XD1E�3�P�E�d�    j�'������E�    �EP�D������te�M�� �M�U�B%��  ��tC�M�yt:�U�B%��  ��t*�M�yt!hHzj h:  h�pj�u�������u̋E�M�H�E������   �j�$����ËM�d�    Y_^[��]�������������������������������������������������������������̋�U��Q�pI�E��M�pI�E���]������������������̋�U��pI]����̋�U��Q�E�   �E�M���M��t �U�E��E���E;�t�E�    �ЋE���]����������������������������̋�U��j�h %h"�d�    P���SVW�XD1E�3�P�E�d�    ��H��u
�   ��  j�S������E�    �����E��}����   �}����   �M��MЋUЃ��UЃ}���   �E��$���h�}h$Uj j j j �X�������u��   h�}h$Uj j j j �3�������u��dh�}h$Uj j j j ��������u��Bhh}h$Uj j j j ���������u�� h4}h$Uj j j j ���������u��E�    ��  �E�   �di�E���M��U�}� ��  �E�   �E�H����  ��t#�U�zt�E�H����  ��t	�U�zu�E�H����  ���o�U���E�(}j��HP�M��Q���������uz�U�z t=�E�HQ�U�BP�M�� Q�U�BP�M�Qhxyj j j j �������(��u��-�E�� P�M�QR�E�Ph�xj j j j ������ ��u��E�    j��HR�E�H�U�D
 P�"�������uz�M�y t=�U�BP�M�QR�E�� P�M�QR�E�Phxj j j j �E�����(��u��-�U�� R�E�HQ�U�Rhhwj j j j ������ ��u��E�    �M�y ��   �U�BP��HQ�U�� R�y�������ud�E�x t2�M�QR�E�HQ�U�� Rhh|j j j j ������ ��u��"�M�� Qh�{j j j j ��������u��E�    �}� uz�E�x t=�M�QR�E�HQ�U�BP�M�� Q�U�Rhp{j j j j �2�����(��u��-�M�QR�E�� P�M�Qh<{j j j j ������ ��u��E�    �G����E������   �j�����ËE܋M�d�    Y_^[��]ÍI ����k�F����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h %h"�d�    P���SVW�XD1E�3�P�E�d�    ��H�E�}�t�M����  ���t	�E�    ��E�   �U܉U��}� u!h8~j hx  h�pj�i�������u̃}� u0�����    j hx  h�ph~h8~�>�������H�sj�h������E�    ��H�M�}�t7�U��t�ti   ��E��%��  �ti�\i    �M��H�E������   �j�&����ËE�M�d�    Y_^[��]������������������������������������������������������������������������������������������̋�U��j�h@%h"�d�    P���SVW�XD1E�3�P�E�d�    3��} ���E��}� u!hD�j h�  h�pj���������u̃}� u+�q���    j h�  h�ph�hD���������s��H��u�fj��������E�    �di�E���M��U�}� t$�E�H����  ��u�UR�E�� P�U�����E������   �j�����ËM�d�    Y_^[��]�������������������������������������������������������������������������������������̋�U��3��} ��]����������������̋�U��Q�} u3��   j j �E�� P�������u3��h�=�wuI�M�� Q�9�����E��}� t�U�� R�E�P������2��M�� Qj ��tR�̒���E�� Pj ��tQ�̒��]��������������������������������������̋�U��j�h`%h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    �E�    �} t	�E�     �} t	�M�    �} t	�U�    �EP��������u3���   j�������E�    �M�� �M��U��B%��  ��t"�M��yt�U��B%��  ��t	�M��yukj�UR�EP�'������tU�M��Q;UuJ�E��H;�H<�} t�U�E��H�
�} t�U�E��H�
�} t�U�E��H�
�E�   ��E�    �E������   �j�����ËE�M�d�    Y_^[��]������������������������������������������������������������������������������������������������̋�U��Q�EP�������u�����M�� �M��U��B��]������������������̋�U��Q�hi�E��M�hi�E���]������������������̋�U��hi]����̋�U��j�h�%h"�d�    P���SVW�XD1E�3�P�E�d�    3��} ���E܃}� u!h �j h�  h�pj�O�������u̃}� u.������    j h�  h�phԀh ��$������m  j�P������E�    �U�di��E�    �	�M���M�}�}�U�E�D�    �M�U�D�    �ӡdi�E���M���U��}� ��   �E��H����  |f�U��B%��  ��}V�M��Q����  �E�L����U��B%��  �U�L��E��H����  �U�D��M�A�U��J����  �U�D��W�E��x t/�M��QR�E��HQ�U�Rh��j j j j ������ ��u���M�Qh`�j j j j ��������u������E�`i�H,�U�Ti�B0�E������   �j�����ËM�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������̋�U���V�E�    3��} ���E�}� u!h �j h;	  h�pj���������u̃}� u0�S����    j h;	  h�pht�h �������3��  3҃} �U��}� u!hL�j h<	  h�pj�h�������u̃}� u0������    j h<	  h�pht�hL��=�����3��0  3Ƀ} ���M�}� u!h$�j h=	  h�pj���������u̃}� u0�����    j h=	  h�pht�h$��������3���   �E�    �	�E����E��}�}�M��U�E��u�L�+L��U��E�L��M��U�E��u�L�+L��U��E�L��M��U�|� u�E��M�|� t$�}� t�}�u�}�u��H��t�E�   �r����E�M�P,+Q,�E�P,�M�U�A0+B0�M�A0�U�    �E�^��]�����������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�P�M��Z����M�����P�MQ�  ���M�������]��������������������̋�U��Q�M��E��@ �} ��   �����M��A�U��B�M��Pl��E��H�U��Ah�B�M��;�Wt�E��H�Qp#�Vu
�����M���U��B;�Tt�M��Q�Bp#�Vu������M��A�U��B�Hp��u�U��B�Hp���U��B�Hp�M��A��U��J�U���J�E���]� ������������������������������������������������������̋�U��Q�M��E��H��t�U��B�Hp����U��B�Hp��]�������������������̋�U��Q�M��E���]����������������̋�U��j�h�%h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    j�������E�    h��h$Uj j j j ���������u̃} t�M��U�di�E���M��U�}� �(  �E�;E��  �M�Q����  ��t)�E�H����  t�U�B%��  ��u��H��u��  �U�z twj j�E�HQ�������tj�U�BP�В��t$�M�QRh��j j j j �*�������u��)�M�QR�E�HQhp�j j j j ���������u̋E�HQhh�j j j j ���������u̋E�H����  ����   �U�BP�M�Q������  R�E�� Ph(�j j j j ������ ��u̃=hi t,j�U�� R�В��u�E�HQ�U�� R�hi����E�P�MQ�  ���   �U�zu;�E�HQ�U�� Rh��j j j j ��������u̋M�Q�UR�x  ���Z�E�H����  ��uI�U�BP�M�Q������  R�E�� Ph��j j j j ������ ��u̋U�R�EP�  ��������E������   �j�B�����h��h$Uj j j j �i�������u̋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���t�XD3ŉE��EP�M�������E�    �	�M����M��U�z}�E�H�M���E�   �U�;U��  �EE��H �M��M��������t3�M����������   ~ �M������PhW  �E�P��������E��hW  �M�Q�M�����P��������E��}� t	�U��U���E�    �E��M��L�������U������     �E�Ph��M�k��1   +�R�E�k��L�Q�������}*j hc	  h�phĂhH^j"j�.����R�&����� �����M��������U��D� �E�P�M�Qh��j j j j ��������u̍M������M�3��������]������������������������������������������������������������������������������������������������������������������̋�U���4�E�P�h�����}� u�}� u��H��t7�}� t1h��h$Uj j j j �-�������u�j �������   �3���]����������������������������������������̋�U���3��} ���E��}� u!h �j h
  h�pj�	�������u̃}� u.�����    j h
  h�ph��h ���������   �E�    �	�U����U��}�}>�E����oQ�U��E�L�Q�U��E�L�Qhh�j j j j �+����� ��u�볋E�H,Qh@�j j j j ��������u̋E�H0Qh�j j j j ���������u̋�]�������������������������������������������������������������������̋�U��j j j �EP�MQ�������]�������������������̋�U��EP�MQj �UR�EP������]���������������̋�U��j j j �EP�MQ�UR������]���������������̋�U��j j j �EP�MQ�UR�EP������]�����������̋�U��EP�MQj �UR�EP�MQ������]�����������̋�U��EP�MQj �UR�EP�MQ�UR�=�����]�����������������������̋�U��j j �EP�MQ�UR������]�����������������̋�U��� �E��#E������E�u!hH�j h9  h�pj�V�������u̃}� u0������    j h9  h�ph�hH��+�����3��$  �} t�U;Ur	�E�    ��E�   �E�E�}� u!h��j h:  h�pj���������u̃}� u0�W����    j h:  h�ph�h��������3��   �}v�U�U���E�   �E����E3�+M���M��UR�EPj�M�M�U�DP�������E�}� u3��M�M�MM��U�D�M��#�+E�E��U�+U����U�j��HP�M���Q��������U��E��E���]��������������������������������������������������������������������������������������������������������������������̋�U��j j �EP�MQ�UR�EP������]�������������̋�U��j j �EP�MQ�UR�EP�MQ������]���������̋�U���,�} u!�EP�MQ�UR�EP�MQ�������  �} u�UR�6�����3��~  �E������E�j��HQ�U��R���������t1�EPh �j j j j�>�������u������    3��$  j��HR�E��P��������u�MQh��j j j j���������u̋E��#E������E�u!hH�j h�  h�pj��������u̃}� u0�����    j h�  h�pht�hH��������3��|  �} t�U;Ur	�E�    ��E�   �E܉E��}� u!h��j h�  h�pj��������u̃}� u0�����    j h�  h�pht�h���d�����3���   �U�P�������M�U++E�}v�E�E���E�   �M؃��M3�+U���U�EP�MQj�U�U�E�LQ�������E��}� u3��   �U�UU�E�L�U��#�+M�M��E�+E���E�j��HQ�U���R�������E��M���U�;Uv�E�E���M�MԋU�R�EP�M�Q�������j�U�P��������E���]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�    �E�    �} vk�����3��u;E����E�u!h�uj h$  h�pj�I�������u̃}� u-������    j h$  h�phX�h�u������3��s�U�U�U��} t�EP�MQ�UR�X������E��E P�MQ�UR�EP�M�Q�UR�x������E�}� t �E�;E�s�M�+M�Qj �U�U�R�������E��]���������������������������������������������������������������������������̋�U��EP������]�������������̋�U��Q�} u�   �E������E�j��HQ�U��R�=�������t!�EPh��j j j j��������u��Lj��HR�E���P���������u�MQh��j j j j�G�������u�j�E��Q��������]�����������������������������������������������������̋�U��Q��H�E��M��H�E���]������������������̋�U��Q�pi�E��E���]�����������̋�U��pi]����̋�U��EP�MQ�UR�E�����]���������������������̋�U��� �E�    �E�    �E�    �E�    �E�    3��} ���E�}� u!h$�j h�  h�pj�f�������u̃}� u.������    j h�  h�ph�h$��;���������w�E�    �U������U��E��Q��������E��U��E+�E�3�+M���M�}v�U�U���E�   �E����E�M�U�D
+E�E�M�+M�+M�M��E���]�������������������������������������������������������������������������th  �   ����t�   �3�������������̋�U��j�h�%h"�d�    P��$SVW�XD1E�3�P�E�d�    �e�3��E��E�  �M�MЍU�UԉE��M�QjPh�m@�|��	�   Ëe��E������E�M�d�    Y_^[��]��������������������������������������̋�U��E��w$���H��l����tRP�EQP�D   ��]úL�R�   P�E�   QP�$   ��]�������������������������������̋�U���<  �XD3ŉE�S�]VW�}S������ǅ����    �u�������������uS�P������������5ܒj j j�Wj h��  ��=   s&P������Pj�Wj h��  �օ�t�������������
ǅ����Њh  �9����}����t%����������RSPW��  �����$  2��������� ������u���  ��t�������   h  ������Q������Rh  ������P���S�`�������t-������������QWh��������R�UP������QR���   �=ؒj j h
  ������Pj�������Qj h��  �h��ׅ�t������j j h
  ������Rj�������Pj h��  �P��ׅ�t�������������U������Q�MRh(�VPSQ����������u�Ԓ�M�_^3�[������]�����������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h�%h"�d�    P��$SVW�XD1E�3�P�E�d�    �e�3��E��E�  �M�MЋU�UԋM�M؍U�U܋M�M��E��U�RjPh�m@�|��	�   Ëe��E������E�M�d�    Y_^[��]����������������������������������������������������̋�U���  �XD3ŉE��=�H��E�������E��   �8 SV��   �ȍq���A��u�+΃�-��   w{������3ɍd$ ����������A��u�Њ@��u�W������+�O�OG��u��������ȃ�����Ȋ@��u�������+���O�OG��u������ȃ��_��T���H������SjPQ������^[�M�3��E�����]��������������������������������������������������������������������̋�U���D  �XD3ŉE�S��HV�uW�}�����������   hȌ������   h��P����i����   ����   �M�Vh��Qh|���$Rhp��~ Wh`�h�������h��Q�ЋV��$RW�E�P�M�Q��   ��8h �U�Rh��E�Ph��������Q���������R��i������������PjSQ�c�����(_^[�M�3��������]�h��jSW�A������M�_^3�[�������]�����������������������������������������������������������������������������̋�U����ESV�u�E��EW3�+ƉE����M��r�   ;�s&�0�U���Qh�R��i�E��E����GF�ɋM�E�y� � _^[��]���������������������������������̋�U���  �XD3ŉE��=�H��E��   SV����   �ȍq�A��u�+΃�:��   ww������3Ɋ�̉������A��u�Њ@��u�W������+�O�OG��u��������ȃ��܉�Ȋ@��u�������+���O�OG��u������ȃ��_��،��HSjP�EP�z�����^[�M�3�������]�����������������������������������������������������������������������̸   ����������̋�U��E��w	���]�3�]������̋�U��M��w�U���H���H]Ã��]�����������̋�U��M��i��i��i    ]�����������������̋�U��M��i��i��i    ]�����������������̡�i����������̡�i�����������u�U��� PRSVWhH�hLjBh��j�߻������u�_^[ZX��]������������������������̋�U�층�]����̋�U���]����̋�U���������   u<�E�8csm�t1�M�9&  �t&�U�%���="�r�M�Q ��t
�   ��   �E�H��ft4�U�z t�} uj��EP�MQ�UR�n������   ��   �   �E�x u$�M��������!���   �E�x ��   �M�9csm�uX�U�zrO�E�x"�vC�M�Q�B�E��}� t1�M$Q�U R�EP�MQ�UR�EP�MQ�UR�U��� �E��E��0�)�E P�MQ�U$R�EP�MQ�UR�EP�MQ�i   �� �   ��]���������������������������������������������������������������������������������������������̋�U���D�E� �E� �E�x�   �M�Q���   �E��	�M�Q�U��E��E��}��|�M�U�;Q}�蜵���E�8csm��[  �M�y�N  �U�z �t�E�x!�t�M�y"��&  �U�z �  �V������    u��  �C������   �E�5������   �M�E�j�UR��������t�������E�8csm�u;�M�yu2�U�z �t�E�x!�t�M�y"�u�U�z u蹴����������    ty�������   �E�����ǀ�       �M�Q�UR��  ������t�C�M�Q�i  ���Ѕ�t+j�EP�,�����hT��M��z���h &�M�Q������������U�:csm��n  �E�x�a  �M�y �t�U�z!�t�E�x"��9  �M�y �+  �U�R�E�P�M�Q�U R�EP�i������E���M����M��U���U�E�;E���   �M�;U��E�M�;H~�ˋU�B�E��M�Q�U���E���E�M����M��}� ��   �U�B�H���M؋U�B�H��U���E܃��E܋M؃��M؃}� ~d�U؋�EԋM�QR�E�P�M�Q��������u���E��U�R�E$P�M Q�U�R�E�P�M�Q�UR�EP�MQ�UR�EP�  ��,�	���D���������M��tj�UR�x������E�����   �M��������!���   �E�x ��   �M�QR�EP�  ���ȅ���   �]������   �U��O������   �E��A����M���   �3����U���   �}$ u�EP�MQ�>�����UR�E$P�/���j��MQ�UR�EP�/������M�QR�  ��������M���   ������U���   �@�E�x v7�M��u*�U$R�E P�M�Q�UR�EP�MQ�UR�EP�  �� ��B����������    u��`�����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�M��EP�M������M��h��E���]� ��������̋�U��Q�M��E�� h��M��������]������������������̋�U��Q�M��M�������E��t�M�Q觴�����E���]� �����������������̋�U��Q�M��EP�M������M��h��E���]� ��������̋�U���V�E�8  �u�X  �U������    tL�G���������9��   t8�M�9MOC�t-�U$R�E P�MQ�UR�EP�MQ�UR� �������t��   �E�x t������M�Q�U�R�EP�M Q�UR�h������E���E����E��M����M��U�;U���   �E��M;|\�U��E;BQ�M��Q�����E��H�| t�U��B�����M��Q�D�H��u�U��B�����M��Q���@t�w���j�M$Q�U R�E�Pj �M��Q�����E�PR�MQ�UR�EP�MQ�UR��  ��,�3���^��]����������������������������������������������������������������������������������������������������������̋�U��Q�E�x t�M�Q�B��u
�   �   �M�U�A;Bt$�M�Q��R�E�H��Q�x�������t3��O�U���t
�M���t1�E���t
�U���t�M���t
�E���t	�E�   ��E�    �E���]����������������������������������������������������̋�U����E��M��U���E��}�MOC�t�}�csm�t�@����ǀ�       �0����n������    ~�`����   �E�M����E�3��3���]������������������������������̋�U��j�hH&h"�d�    P���SVW�XD1E�3�P�E�d�    �e�E�x�   �M�Q���   �E��	�M�Q�U܋E܉E������   �E؋M؋���E؉�E�    �M�;M��   �}��~�U�E�;B}��j����M�Q�E�M��E�   �U�B�M�|� t%�U�E��Bh  �MQ�U�B�M�T�R肱���E�    ��E�P������Ëe��E�    �M��M��f����E������   �)��������    ~������   �EԋUԋ���MԉËU�;Uu�讪���E�M�H�M�d�    Y_^[��]������������������������������������������������������������������������������������������������̋�U����E�E��}  t�M Q�UR�E�P�MQ�������}, u�UR�EP�+�����MQ�U,R�����E$�Q�UR�EP�M�Q�������U$�B���M�Ah   �U(R�E�HQ�UR�EP�M�Q�UR�T   ���E��}� t�EP�M�Q�.�����]�������������������������������������������������������̋�U��j�hx&h"�d�    P���SVW�XD1E�3�P�E�d�    �e�E�E��E�    �M�Q��U��E�HQ�U�R�������E���������   �E���������   �M�������U���   ������M���   �E�    �E�   �E�   �U R�EP�MQ�UR�EP�������E��E�    ��   �M�Q�N  ��Ëe��e���ǀ      �U�B�E��M�y�   �U�B%�   �ȉM��	�U�B�E��M��M��U�B�E��E�    �	�Mă��MċU�E�;BsG�M�k��U��E�;D
~3�M�k��U��E�;D
!�M�k��U��D
���E��M��U��ʉE��륋M�Q�URj �EP�ޭ�����E�    �E�    �E������E�    �   �   �M�U��Q��E�P膶�����a����Mȉ��   �S����Ủ��   �E�8csm�u\�M�yuS�U�z �t�E�x!�t�M�y"�u/�}� u)�}� t#�U�BP��������t�M�Q�UR������ËEЋM�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E��M��U��:csm�uN�E��xuE�M��y �t�U��z!�t�E��x"�u!�M��y u�����ǀ     �   ��3���]�����������������������������������̋�U��j�h�&h"�d�    P���SVW�XD1E�3�P�E�d�    �e��E�    �E�x t#�M�Q�B��t�M�y u�U�%   �u3���  �M���   �t�E�E���M�Q�E�L�M��E�    �U���tXj�M�QR�R�������t9j�E�P��������t'�M��U�B��M��Q�U��P�������M���苤���@  �U���txj�M�QR���������tYj�E�P�+�������tG�M�QR�E�HQ�U�R�}������E�xu"�M��9 t�U��R�E��Q�������U����	����   �E�x uZj�M�QR�o�������t>j�E�P��������t,�M�QR�E��P�M�QR������P�E�P�������裣���[j�M�QR��������tAj�E�P�P�������t/�M�QR豺������t�E���t	�E�   ��E�   ��F����E�������   Ëe�������E������E�M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h�&h"�d�    P���SVW�XD1E�3�P�E�d�    �e�E���   �t�U�U���E�H�U�D
�E��E�    �MQ�UR�EP�MQ菺�����E��}�t�}�t+�R�U��R�E�HQ�������P�U�BP�M�Q�0����)j�U��R�E�HQ������P�U�BP�M�Q�x����E�������   Ëe��M����E������M�d�    Y_^[��]��������������������������������������������������������������������̋�U��j�h�&h"�d�    P��SVW�XD1E�3�P�E�d�    �e�} t�E�8csm�t�U�M�y tL�U�B�x t@�E�    �M�Q�BP�M�QR������E�������E�����Ëe��Z����E������M�d�    Y_^[��]�������������������������������������������������̋�U��Q�E�M�M��U�z |'�E�H�U�
�M�Q�M��M��U�E�B�E��E���]������������������������̋�U�������3Ƀ��    ����]������̋�U���(�} u3���  �E��M��} t�U�B����   �M��9MOC�t�U��@uz�E��8csm�uK�M��yuB�U��z �t�E��x!�t�M��y"�u�U��z u�H������    u3��H  �3����   �E܋E܋���U܉
�   �$  �E��8csm��  �M��y�  �U��z �t�E��x!�t�M��y"���   �U��z u#��������    u3���   �������   �E��M�M�U�U��E�   ��E��M��Q�B���E�M��Q�B��M���U����U��E���E�}� ~d�M��U��E��HQ�U�R�E�P�Ʊ������t?�.����   �E؋M؋���E؉�} t�M�Q�U�R�EP�M�Q�g������   ��3���]�������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�E��M����M�U���U��} ��   �E�8 ��   �M��U��E��8csm�uD�M��yu;�U��z �t�E��x!�t�M��y"�u�U��z u��������   �E��M��QR�E�P�������E�������M􋐈   ������M����   ������M����   ��U�������E�� ���������   �E�M����E��h������    }�Z���ǀ�       �   ��]������������������������������������������������������������������������������������̋�U����} u3��l�E��M��U��:csm�uW�E��xuN�M��y �t�U��z!�t�E��x"�u*�M��y u!�����   �E��U�����M���   �3���]����������������������������������������������̋�U����E�E��M����M�U���U��E�8��G  �M�Q�+������} ��   ��������   �:csm�u~��������   �xum��������   �y �t(��������   �z!�t�������   �x"�u1�������   �QR�&�������tj�������   P�8������k������   �9csm�um�X������   �zu\�G������   �x �t(�3������   �y!�t�������   �z"�u �} t�����   �E��E�����U��
������M����   ������M�����   ��]���������������������������������������������������������������������������������������������������������̋�U��   ]����̋�U��j�h'h"�d�    P��SVW�XD1E�3�P�E�d�    �e��E�    �M�U�E�������E�P臰����Ëe��E������M�d�    Y_^[��]��������������������������������������������̋�U��j�h('h"�d�    P��SVW�XD1E�3�P�E�d�    �e��E�    �EP�U���E�������M�Q������Ëe��E������M�d�    Y_^[��]����������������������������������������̋�U��j�hH'h"�d�    P��SVW�XD1E�3�P�E�d�    �e��E�    �EP�U�E�������M�Q�F�����Ëe��E������M�d�    Y_^[��]�������������������������������������������̋�U��j�hh'h"�d�    P��SVW�XD1E�3�P�E�d�    �e��E�    �EP�MQ�UR�EP�U�E�������M�Q蚮����Ëe��E������M�d�    Y_^[��]�����������������������������������������������̋�U����} t�螖���} u�`����E� �E�    �	�E���E�M�U�;}m�E�H�Q���U��E�H�Q��E���M����M��U����U��}� ~4�E���M�U�BP�M�Q�U����EPR賩������t�E���뀊E��]������������������������������������������������������������̋�U��j�hp�d�    PQSVW�XD3�P�E�d�    �e��������    u�胕���E�    躝���$�����M���   j j ������E������y���E����������M�d�    Y_^[��]������������������������������������������������̋�U��Q�E�    �	�E����E��M�U�;}'h�H�E����M�Q�L�̲������t����2���]���������������������������������̋�U����} t��~����E��M�}� t��i����U�:csm�u/�E�xu&�M�y �t�U�z!�t�E�x"�u��*����M�Q�B���E��M�Q�B��M���U����U��E����E��}� ~0�M���U��E��H��Q�M蟪��P��������u�   ��3���]�����������������������������������������������������������U���SQ�E���E��EU�u�M�m��$���VW��_^��]�MU���   u�   Q����]Y[�� �������������������̋�U����E�    �4IP����t(�=0I�t�0IQ�4IR���ЉE��}� u*h����������E�}� tht��E�P���E���M����  �U��}� t
�EP�U��E�E��]��������������������������������������������̋�U��Q�EP���E��}� t�E���MQ�i�������]������������������̋�U��j �~�����]���������������̋�U����E�    �4IP����t(�=0I�t�0IQ�4IR���ЉE��}� u*h����������E�}� th���E�P���E���M����  �U��}� t
�EP�U��E�E��]��������������������������������������������̋�U�����]� ����������������̋�U��EP�4IQ����]� �������������������̋�U��0I]����̋�U��Q�4IP���E��}� u"��iQ谦�����E��U�R�4IP����E���]����������������������������̋�U��EP�MQ��iR�^�������]� �������������̋�U���h���l������E��}� u�����3���  h��E�P����ih��M�Q����ih���U�R����ih���E�P����i�=�i t�=�i t�=�i t	�=�i u,��ij�����i�����i�����i����4I�=4I�t��iQ�4IR�����u3��	  �������iP譖������i��iQ虖������i��iR腖������i��iP�r�������i苧����u����3��   h>���iQ�Ѥ�����У0I�=0I�u	����3��th�  h��jh  j�$������E��}� t�U�R�0IP��iQ�{������Ѕ�u	�B���3��(j �U�R�\������Ē�M���U��B�����   ��]��������������������������������������������������������������������������������������������������������������������������������������̋�U��=0I�t!�0IP��iQ藣�������0I�����=4I�t�4IR����4I�����M���]��������������������������̋�U��j�h�'h"�d�    P���SVW�XD1E�3�P�E�d�    h���B������E�E�@\�B�M�A   �}� t0ht��U�R���M���  h���U�R���M���  �U�Bp   �Eƀ�   C�MƁK  C�U�Bh�Pj�%������E�    �E�HhQ�X��E������   �j�������j�������E�   �U�E�Bl�M�yl u�U��W�Bl�M�QlR�������E������   �j�������ËM�d�    Y_^[��]���������������������������������������������������������������������������������������������̋�U�������E��0IP蚇���ЉE��}� uj hL  h��jh  j��������E��}� tY�M�Q�0IR��iP�4������Ѕ�t%j �M�Q�������Ē�U���E��@�����j�M�Q�ݛ�����E�    �U�R� ��E���]���������������������������������������������������������̋�U��Q�����E��}� u
j�K������E���]�����������̋�U��j�h(h"�d�    P���SVW�XD1E�3�P�E�d�    �E�E܃}� ��  �M܃y$ tj�U܋B$P� ������M܃y, tj�U܋B,P�������M܃y4 tj�U܋B4P�̚�����M܃y< tj�U܋B<P貚�����M܃y@ tj�U܋B@P蘚�����M܃yD tj�U܋BDP�~������M܃yH tj�U܋BHP�d������M܁y\�Btj�U܋B\P�G�����j�������E�    �M܋Qh�U��}� t%�E�P�\���u�}��Ptj�M�Q�������E������   �j��������j薍�����E�   �U܋Bl�E�}� t4�M�Q��������U�;�Wt�}�Vt�E�8 u�M�Q�d������E������   �j�W������j�U�R�n������M�d�    Y_^[��]� ���������������������������������������������������������������������������������������������������������������������������������������������̋�U��=0I�tQ�} u)�4IP����t�0IQ�4IR���ЉEj �0IP��iQ薝�����ЋUR�����=4I�tj �4IP���]����������������������������������������̋�U���Ē]���̋�U����]���̋�U��h��苎������i]�������̋�U��j�hH(h"�d�    P���SVW�XD1E�3�P�E�d�    �e������@x�E�}� t#�E�    �U��E�������   Ëe��E������$����M�d�    Y_^[��]��������������������������������̋�U��Q�x����@|�E��}� t�U��!�����]�������������̋�U��j�hh(h"�d�    P���SVW�XD1E�3�P�E�d�    �e衤iP��������E�}� t#�E�    �U��E�������   Ëe��E�����蜋���M�d�    Y_^[��]������������������������������������������̋�U���(  ��j��j��j��j�5�j�=�jf��jf��jf��jf��jf�%�jf�-�j���j�E ��j�E��j�E��j������� j  ��j��i��i	 ���i   �XD�������\D�����������ij蒎����j ���h(�����=�i u
j�l�����h	 ����P�����]����������������������������������������������������������������������������������̋�U��j jh�h��h8�h   h   j 誘����P������]�������������������������̋�U����x��]��h��]��E��u��M��m��]����]�����z	�E�   ��E�    �E��]��������������������̋�U���h�����E��}� t!h���E�P���E��}� t	j �U���茍����]��������������������������̋�U��j �EP�Н����]�����������̋�U����EP�M��A����M�R�Ŗ������et�E���E�M�R薅������u�E�Q蕖������xu	�U���U�E��M��M��N�������   ��U���M���M�U��E��M�U���E��E��M��E���E��u׍M��������]������������������������������������������������̋�U��j �EP�I�����]�����������̋�U���V�EP�M��0����M���t*�E�0�M�肄������   ��;�t�U���U�̋E��U���U����   �E���t!�U���et�M���Et�E���E�ՋM�M��U���U�E���0u�U���U��E�0�M���������   ��;�u	�U���U�E���E�M�U����M��E����E���t�؍M�蛣��^��]�������������������������������������������������������������������̋�U��Q�E�������Az	�E�   ��E�    �E���]���������������������̋�U����} t$�EP�MQ�U�R�7������E�M���U��P��EP�MQ�U�R�ٷ�����E�M���]������������������������������̋�U��j �EP�MQ�UR�3�����]�������������������̋�U���D�XD3ŉE��E�E܍M̉M��E�    j�U�R�E�P�M܋QR�P������3Ƀ} ���Mă}� u!ht�j h�  h�j蠂������u̃}� u3�"����    j h�  h�hؑht��u������   �  3�;E��ىM�u!h��j h�  h�j�8�������u̃}� u3躠���    j h�  h�hؑh���������   �   �}�u�E�E���M�3҃9-�E+�3Ƀ} ��+��E��U�R�E��P�M�Q�U�3��:-��E3Ƀ} ���P�ޣ�����Eȃ}� t�U� �E��(�EPj �M�Q�UR�EP�MQ�UR�   ���EȋEȋM�3��դ����]��������������������������������������������������������������������������������������������������������������������̋�U���@�E�    �E P�M��ʊ��3Ƀ} ���M܃}� u!ht�j hL  h�j薀������u̃}� u@�����    j hL  h�h��ht��k������E�   �M�跟���E���  3�;E��ىM�u!h��j hM  h�j�!�������u̃}� u@裞���    j hM  h�h��h����������E�   �M��B����E��}  3��} ����#E��	;E��ىM�u!hp�j hU  h�j�������u̃}� u@����� "   j hU  h�h��hp��q������E�"   �M�轞���E���  �E��t'�M3҃9-��U�U�3��} ��P�M�Q�V  ���U�U��E�8-u�M��-�U����U��} ~-�E��M��Q��E����E��M��S~������   ��M����E�E�M��Ƀ���E��}�u�U�U���E�+E�M+ȉM�j h�  h�h��h��h���U�R�E�P蚞����P�)������M����M�} t�U��E�E����E��M�Q���0��   �M�Q���U�y�E��؉E��M��-�U����U��}�d|)�E���d   ���ЋE��ʋU��
�E���d   ���U��U����U��}�
|)�E���
   ���ЋE��ʋU��
�E���
   ���U��U����U��E��M��ЋE���Lu��t �U����0uj�M��Q�U�R�a������E�    �M�������Eċ�]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�t����]�����������̋�U���   �E�E��E��  �E�    �E�    �E�    �0   f�M��E�    �E�    3�f�U��E�    �E�    �E�    �E�    �EP�M��Ӆ���} }�E    3Ƀ} ���M��}� u!ht�j h&  h�j�{������u̃}� u@�����    j h&  h�h|�ht��g������E�   �M�賚���E���  3�;E��ىM�u!h��j h'  h�j�{������u̃}� u@蟙���    j h'  h�h|�h���������E�   �M��>����E��g  �E�  �M��;M��ډU�u!h�j h/  h�j�z������u̃}� u@� ���� "   j h/  h�h|�h��s������E�"   �M�这���E���  �M��Q�4�I���%�  �� �E��U��}��  ��   �}� ��   �}�u�U�U��	�E���E�j �MQ�U�R�E��P�MQ襂�����E��}� t�U� �E��E��M��2����E��[  �M�Q��-u�E� -�M���M�U�0�E���E�M��ɀ����x�U�
�E���Eje�MQ�"������E��}� t!�U��Ҁ����p�E���M����M��U�� �E��E��M�蟘���E���  �M��Q�?�)������� ��|����U���|���U�t�E� -�M���M�U�0�E���E�M��ɀ����x�U�
�E���E�M��ɀ����a�у�:�U��M��Q�4豗��%�  �� ��t�����x�����t����x���u[�E� 0�M���M�U��J���� ��l�����p�����l����p���u�E�    �E�    ��EЃ��Mԃ� �EЉM���U�1�E���E�M�M��U���U�} u�E��  ��M��kw������   ��M����E��P���� ��d�����h�����h��� w��d��� �p  �E�   �E�    �M܋E�U��|v���E�U��E܅���   �} ~}�M��Q���� #E�#U��M��m���f�E��U���0f�U��E���9~�M�M�f�M��U�E���M���M�E�U��,����E�U��U܃�f�U܋E���E�q����M܅���   �U��R���� #E�#U��M�����f�E��E�����   �M�M��U����U��E����ft�U����Fu�M��0�U����U��ًE�;E�t/�M����9u�E���U��D�M����U�����M����U����U��E�����U��
�	�E���E�} ~�M�0�U���U���E����u�U��U�E���$�p�M��U���U�M��Q�4�����%�  �� +E�UԉE��U�}� |�}� r�U�+�E���E�"�M�-�U���U�E��؋M�� �ىE��M�U�U��E�� 0�}� |M	�}��  rBj h�  �M�Q�U�R�u������0�M��U���Uj h�  �E�P�M�Q�Wu���E��U�U;U�u�}� |D�}�dr<j jd�E�P�M�Q�\u���Ѓ�0�E��M���Mj jd�U�R�E�P�u���E��U�M;M�u�}� |D�}�
r<j j
�U�R�E�P�
u���ȃ�0�U�
�E���Ej j
�M�Q�U�R�t���E��U��E���0�M��U���U�E�  �E�    �M��ғ���E���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EP�MQ��i����]���������̋�U��j �EP�MQ�UR�EP�MQ�3j����]�����������̋�U���D�XD3ŉE��E�E܍M̉M��E�    j�U�R�E�P�M܋QR�P�������3Ƀ} ���Mă}� u!ht�j h�  h�j�q������u̃}� u3�2����    j h�  h�h��ht�腅�����   ��   3�;E��ىM�u!h��j h�  h�j�Hq������u̃}� u3�ʏ���    j h�  h�h��h���������   �   �}�u�E�E���M�3҃9-�E+E��M�Q�U��EBP�M�Q�U�3��:-��EP�������Eȃ}� t�M� �E��$�URj �E�P�MQ�UR�EP�   ���EȋEȋM�3��������]�����������������������������������������������������������������������������������������������������������̋�U���4�E�H���M��UR�M���y��3��} ���E�}� u!ht�j h  h�j��o������u̃}� u@�C����    j h  h�h��ht�薃�����E�   �M������E��  3�;U��؉E�u!h��j h  h�j�Lo������u̃}� u@�΍���    j h  h�h��h���!������E�   �M��m����E��B  �U��t7�E3Ƀ8-��M�M��U�;Uu�E�E��E܋M��0�U܃��U܋E��  �M�M��U�:-u�E�� -�M����M��U�z j�E�P��  ���M��0�U����U���E�M�H�M��} ��   j�U�R�  ���M���m��� ���   ��E��
��U����U��E�x }]�M��t�U�B�؉E�&�M�Q��9U}�E�E���M�Q�ډŰẺE�MQ�U�R�  ���EPj0�M�Q�ɗ�����E�    �M��&����EЋ�]������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�T�����]���������������̋�U���P�XD3ŉE��E�    �E�E��E� �MȉM�j�U�R�E�P�MċQR�P�������3Ƀ} ���M��}� u!ht�j h�  h�j�|l������u̃}� u3������    j h�  h�hĔht��Q������   �i  3�;E��ىM�u!h��j h�  h�j�l������u̃}� u3薊���    j h�  h�hĔh���������   �  �E؋H���M܋U�3��:-��E�E��}�u�M�M���U�3��:-���M+ȉM��U�R�EP�M�Q�U�R��������E��}� t�E�  �E��   �M؋Q��9U����E��M؋Q���U܃}��|�E�;E|&�MQj�U�R�EP�MQ�UR�EP�?������D�B�M���t�U���M����M���t��U��B� �EPj�M�Q�UR�EP�MQ��������M�3��I�����]��������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�n�����]�����������̋�U��Q�E�    �}et�}Eu%�E P�MQ�UR�EP�MQ�UR�b�����E��{�}fu!�E P�MQ�UR�EP�MQ�������E��T�}at�}Au%�U R�EP�MQ�UR�EP�MQ�ua�����E��#�U R�EP�MQ�UR�EP�MQ諈�����E��E���]������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�UR������]�����������������������̋�U��} t#�EP耕������P�MQ�UUR�q����]����������������̋�U��Q�E�    �	�E����E��}�
s�M���<IR�|l�����M���<I�ҋ�]�������������������������������̋�U��j�h�(h"�d�    P���SVW�XD1E�3�P�E�d�    j�7i�����E�    �E�x ��   �pm�M��E�lm��U��U�}� tV�E�M�;Qu�E��M�Q�P�E�P�Ą�����/�M�M��U�z uhp�j jXh��j�rg������u�랋M�QR脄�����E�@    �E������   �j衟����ËM�d�    Y_^[��]������������������������������������������������������������������������̋�U��j�h�(h"�d�    P���SVW�XD1E�3�P�E�d�    �E�x �I  h (  h��hްj �M��	Qj �N������E�}� u3��  �U�R�*������E��E��M����M���v�U�U���� u�M�M�� ��j�pg�����E�    �U�z ��   j�ے�����E܃}� ��   �E���P迒�����M�A�U�z t[j h�   h��hX�h���E�P�M���Q�U�BP�؅����P�gp�����M܋U�B��M܋U�B�A�M�U܉Q��E�P褂�����M�Q�<������E������   �j违����ËU�B�M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������̋�U��j�h�(h"�d�    P���SVW�XD1E�3�P�E�d�    j��e�����E�    �E�x ��   �pm�M��E�lm��U��U�}� tY�E�M�;Qu�E��M�Q�P�E�P�������2�M�M��U�z u!hp�j h�   h��j�d������u�뛋M�QR�ś�����E�@    �E������   �j�>�����ËM�d�    Y_^[��]���������������������������������������������������������������������̋�U���E��u	� (  f�M�URh��hް�EP�MQ�UR������]���������������������̋�U��j�h�(h"�d�    P���SVW�XD1E�3�P�E�d�    �E�x �a  j�*d�����E�    �M�y �*  h (  j �U��	Rj �P]�����E�}� u"�E�    j��E�PhXD�d�����E��  �M�Q�K������E��U��E����E���v�M�M���� u�E�E��  ��j�������E܃}� ��   �E�    �M���Q��������E؃}� taj h4  h��h�h���U�R�E���P�M�Q������P�l�����U�E؉B�M܋U�B��M܋U�B�A�M�U܉Q��E�P耙�����M�Q�t������E������   �j�������ËU�B�M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������̋�U��j�h)h"�d�    P���SVW�XD1E�3�P�E�d�    j�b�����E�    �E�H�M��E�    ��U��U�}� t%�E�H�M��U�P�S������M�Q�G��������E������   �j�Ș����ËM�d�    Y_^[��]�����������������������������������������������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t�������������������������������������������̋�U���S�E�    �E�    �E�    S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�%   t�1   ��t�   �3�[��]�������������������������������̋�U��j�h()h"�d�    P���SVW�XD1E�3�P�E�d�    �e��E�    �E�    f(��E�   �E������A�E���U��}�  �t�}�  �t	�E�    ��E�   �E�Ëe��E�    �E������E�M�d�    Y_^[��]���������������������������������������������������̋�U���I[���Py3�]�������������̋�U���(�} t�} v	�E�   ��E�    �E�E�}� uh��j jh�j�]������u̃}� u0�|���    j jh�h �h���nq�����   �L  �} ��   �U� �}�tI�}���t@�}v:�E��9�Hs��H�M��	�U���U�E�Ph�   �M��Q������3҃} �U��}� uhЗj jh�j��\������u̃}� u0�S{���    j jh�h �hЗ�p�����   �  �M�M��U�U��E��M���E���U����U��E���E��t�M����M�t�̓}� ��   �U� �}�tI�}���t@�}v:�E��9�Hs��H�M��	�U���U��E�Ph�   �M��Q������������t3�t	�E�   ��E�    �M܉M�}� uhX�j jh�j�[������u̃}� u-�8z��� "   j jh�h �hX��o�����"   �o�}�tg�}���t^�E+E���;EsP�M+M����U+�9�Hs
��H�E���M+M����U+щU؋E�Ph�   �M+M��U�D
P�	�����3���]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��   ]����̋�U���Dy    ]���������������̋�U����E�    �E�    �	�E����E��}�$}\�M��<�|IuM�U�k���xm�E���xI�M����M�h�  �U���xIP��������u�M���xI    3��땸   ��]������������������������������������̋�U����E�    �	�E����E��}�$}O�M��<�xI t@�U��<�|It3�E���xI�M��U�R�l�j�E�P�f�����M���xI    ��E�    �	�U����U��}�$}3�E��<�xI t$�M��<�|Iu�U���xI�E�M�Q�l�뾋�]��������������������������������������������������̋�U��j�hH)h"�d�    P���SVW�XD1E�3�P�E�d�    �E�   �=�t u��m��j躄����h�   芄�����E�<�xI t
�   �   h  h��jj��Q�����E�}� u�xv���    3��   j
�Y�����E�    �M�<�xI uFh�  �U�R�������u"j�E�P�%e�����%v���    �E�    ��M�U��xI�j�E�P��d�����E������   �j
趏����ËE��M�d�    Y_^[��]������������������������������������������������������������������������������������������̋�U��E�<�xI u�MQ�R������u
j�n�����U��xIP�p�]�����������������̋�U��E��xIQ�t�]��������̋�U��EPj ��h�   躂����]����������������̋�U���Ԓ]���̋�U����} |�}}	�E�   ��E�    �E��E��}� u"h�j jthp�j��U������u�6N���}� u.�dt���    j jthp�h@�h��i��������   �}�t�U���t	�E�    ��E�   �E�E�}� u"h8�j jyhp�j�fU������u�M���}� u+��s���    j jyhp�h@�h8��:i��������/�}�u�U���J��E���J�M��U�E���J�E���]������������������������������������������������������������������������������������������̋�U����} |�}}	�E�   ��E�    �E�E��}� u%h�j h�   hp�j�ST������u�L���}� u0��r���    j h�   hp�hH�h��$h����������c�}�u�U���J�Q�E���J�M��}�uj����U���J�'�}�uj����M���J��U�E���J�E���]��������������������������������������������������������������̋�U��Q�,y�E��M�,y�E���]������������������̋�U��,y]����̋�U��j�hh)h"�d�    P���PP  �R���XD1E�3ŉE�SVWP�E�d�    ǅ����    ǅ����    ƅп�� h�  j ��ѿ��P�|����ƅ���� h�  j ������Q�|����3�f������h�  j ������P�{|����ƅЯ�� h�  j ��ѯ��Q�^|�����} |�}|����*  �E�    �}��   h�J�X�����   j h  hp�h��h8�j
h   ��п��R�EP�Zh����P�\����h����} t�M�������
ǅ������������R��h�����п��P��h ����I��ǅ���������=  �} ��   ǅ̯��    �p�����ȯ����o���     �UR�EPh�  h   ��Я��Q�#k������̯����̯�� }*j h-  hp�h��hH^j"j�o���R�L���� �o����ȯ�����̯�� }8j h0  hp�h��h0�h��h   ��Я��R��p����P�t[�����}uV�} tǅ������
ǅ����̠j h5  hp�h��h �������Ph   ��п��Q�p����P�[����j h7  hp�h��h����Я��Rh   ��п��P�sG����P��Z�����}u�M���J��t8j h<  hp�h��h8�h0�h   ��п��P�&G����P�Z����j h=  hp�h��h؞h h   ��п��Q��F����P�YZ�����} ��   ǅį��    �n����������n���     ��п��P�MQ�URhĞh�  h   ������P�a{������į����į�� }*j hD  hp�h��hH^j"j�m���Q�J���� �m�����������į�� }8j hG  hp�h��h�h��h   ������P��n����P�yY�����:j hK  hp�h��h����п��Qh   ������R�n����P�=Y����ǅ����    ǅ����    j�������Ph   ������Q������R�]����������j hP  hp�h��h��j"j������P�I���� ������ t8j hR  hp�h��h�hx�h   ������Q�um����P�X�����=@y u�=<y �#  ǅ����    ǅ����    j��N�����E�   �@y��������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���tǅ����   �������������렃����� un�<y��������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���tǅ����   ���������������E�    �   �j������Ã����� �D  �=,y t?ǅ����    ������R������P�MQ�,y����tǅ����   ������������������ ��   �E���J��t>�U�<��J�t1j ������P������Q��x����P������R�E���JQ���U���J��t������Q���U���J��twƅп�� �} t9j h�  hp�h��h8�j
h   ��п��Q�UR��a����P�<V������Я��P�MQ�U��ҍ�п��#�R�MQ�UR��n�����������E������   ��}uh�J�\�Ë������M�d�    Y_^[�M�3��n����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h�)h"�d�    P���\�  ��G���XD1E�3ŉE�SVWP�E�d�    ǅ����    ǅ����    3�f��Я��h�  j ��ү��Q�r����3�f������h�  j ������P�fr����ƅ���� h�  j ������Q�Ir����3�f��Џ��h�  j ��ҏ��P�*r�����} |�}|����.  �E�    �}��   h�J�X�����   j h�  hp�h�h��j
h   ��Я��Q�UR膀����P�~R����h �� ��} t�E������
ǅ����������Q� �h�� ���Я��R� �h�� ��?��ǅ���������A  �} ��   ��e��� ��ȏ����e���     �MQ�URh�  h   ��Џ��P��Z������̏����̏�� }*j h  hp�h�hH^j"j�xe���Q�pB���� �he����ȏ�����̏�� }8j h	  hp�h�h(�h(]h   ��Џ��P�*f����P�JQ�����}uV�} tǅ������
ǅ���ȧj h  hp�h�h�������Qh   ��Я��R��e����P��P����j h  hp�h�h����Џ��Ph   ��Я��Q�D=����P�P�����}u�U���J��t8j h  hp�h�h0�h(�h   ��Я��Q��<����P�gP����j h  hp�h�hХh�h   ��Я��R�<����P�/P�����} ��   ǅď��    ��c��� ��������c���     ��Я��Q�UR�EPh��h   h   ������Q�k������ď����ď�� }*j h  hp�h�hH^j"j�}c���R�u@���� �mc�����������ď�� }8j h!  hp�h�h�]h(]h   ������R�/d����P�OO�����:j h%  hp�h�hH���Я��Ph   ������Q��c����P�O����ǅ����    j h+  hp�h�h��j"jj�������Rh   ������Pj �Of����P�?���� ������������ t8j h-  hp�h�h��h`�h   ������Q��c����P�N�����=@y u�=<y �#  ǅ����    ǅ����    j��D�����E�   �@y��������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���t������������ǅ����   �렃����� un�<y��������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���t������������ǅ����   ���E�    �   �j��z����Ã����� �g  �=,y t?ǅ����    ������R������P�MQ�,y����t������������ǅ����   ������ �  �E���J���[  �U�<��J��J  �E���JQ�������������t�Jj ������R������P�n����P������Q�U���JP����t��   �����t��   ǅ���    j h~  hp�h�h��j"jj�������Qh   �����R�����P�c����P��<���� ���������� t>�����Pt5j ������Q������R�bm������P������P�M���JR���@����� v������������j ������Q�����R�����P�M���JR���E���J��t������R� ��E���J��ty3�f��Я���} t9j h�  hp�h�h��j
h   ��Я��P�MQ�y����P�K������Џ��R�EP�M��ɍ�Я��#�Q�EP�MQ�[d�����������E������   ��}uh�J�\�Ë������M�d�    Y_^[�M�3��Vc����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��V�D���M��UR��o��������[���0^]������������������������̋�U��Q�E�    �	�E����E��}�-s�M��U;��Ju�E����J�7�ԃ}r�}$w	�   �"� �}�   r�}�   w	�   ���   ��]��������������������������������������������̋�U��Q�7���E��}� u	�   ���[���M�3���]�������������������̋�U��Q3��} ���E��}� u!h��j h�   h(�j�+<������u̃}� u%j h�   h(�h�h���P�����   ��Z���U� �3���]������������������������������������������̋�U��Q��6���E��}� u	�   ���8B���M�3���]�������������������̋�U��Q3��} ���E��}� u!h��j h�   h(�j�K;������u̃}� u%j h�   h(�h��h���+O�����   ��A���U� �3���]������������������������������������������̋�U��Q��5���E��}� u	�`L���E�����]���������̋�U��Q�5���E��}� u	�dL���E�����]���������̋�U���0�E� �E�   �E���E��M����M�U��B3XD�EԋM�Q�U�R��  ���E�H��f�  �U�U��E�E��M��U��Q�E��H�M���U�U؃}����   �E�k��MԍT�U�E�H�MЋU��E�}� ��   �U�M��de���E��E��}� }�E�    �   �   �}� ��   �M�9csm�u)�=P� t hP��oP������tj�UR�P����M����=C���E��H;M�thXD�U�R�M����U��8?���E��M�H�U�R�E�P��   ���U�M�I�[�������&�U��z�thXD�E�P�M����������>���E��M߅�t�U�R�E�P�   ���E��]���������������������������������������������������������������������������������������������������������������������������̋�U����E�8�t%�M��E��M��U�EB3E��E��M��[���M�Q�E��M��U�EB3E��E��M��r[����]���������������������������������̋�U����E��  �E�    �}� u0�E�P�`��MQ���E��U����  �U��}�`�  v��ʋE���]�����������������������������̋�U��Q�=�Y th�Y�5N������t�EP��Y���C��h8h�2V�����E��}� t�E��Gh���`����hh ��  ���=(y th(y��M������tj jj �(y3���]���������������������������������������������������̋�U��j j �EP�^  ��]���������̋�U��j j�EP�>  ��]���������̋�U��jj j �   ��]�����������̋�U��jjj �   ��]�����������̋�U��Q�K���EP�b������LQ�H�����E�h�   �U�����]������������������������̋�U��Q�@o�E��	�M����M��}� t�U��: tj�E��Q�C������j�@oR�C�����@o    �8o�E��	�M����M��}� t�U��: tj�E��Q��B������j�8oR�B�����8o    j�4oP�B����j�0oQ�B����j� yR�G����P�oB�����4o    �0o    �cd��� y��TP�\���u'�=�T�Ptj��TQ�$B������T�P��TR�X���]���������������������������������������������������������������������������������������������̋�U��j�h�)h"�d�    P���SVW�XD1E�3�P�E�d�    ��C���E�    �=Xo�_  �To   �E�Po�} �  � yQ�TF�����E�}� ��   �yR�8F�����E��E�    �E�EԋM؉M�   ����   �E�    �E�    �E؃��E؋M�;M�r��b���U�9u��E�;E�s�n�M؋R��E�����E��b���M؉�U܋ yR�E�����EСyP�E�����E̋M�;M�u�U�;U�t�EЉEԋMԉM�ỦU��E��E��N���hPh<�  ��hXhT�u  ���=\o u#j��2[������ t�\o   �5U���j���E������   ��} t��U��Ã} t��Xo   �U���MQ�^�����M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������̋�U���h�����E��}� th��E�P���E��}� t�MQ�U���]�����������������̋�U��EP��U�����MQ�$�]�������������������̋�U��j�T2����]���������������̋�U��j�Wi����]���������������̋�U��Q�n`���E��E�P�*R�����M�Q�+�����U�R�KK�����E�P��9�����M�Q��(�����U�R�\�����E�P�0�����M�Q�c����hۋ�4������L��]��������������������������������������������̋�U��E;Es�M�9 t�U��ЋM���M��]�����������������������̋�U��Q�E�    �E;Es#�}� u�M�9 t
�U��ЉE��M���M�ՋE���]�����������������̋�U���3��} ���E��}� u!h��j h�  h`�j�i/������u̃}� u0��M���    j h�  h`�h<�h���>C�����   �y3҃=Lo �U��}� u!h�j h�  h`�j��.������u̃}� u0�M���    j h�  h`�h<�h���B�����   ��M�Lo�3���]������������������������������������������������������������������̋�U���3��} ���E��}� u!h��j h�  h`�j�9.������u̃}� u0�L���    j h�  h`�h �h���B�����   �y3҃=Ho �U��}� u!hثj h�  h`�j��-������u̃}� u0�OL���    j h�  h`�h �hث�A�����   ��M�Ho�3���]������������������������������������������������������������������̋�U��E�lo�M�po�U�to�E�xo]�����������������������̋�U��j�h�)h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    �E�    �}t�}u�a  �}t�}t�}t�}t
�}�V  j ��-�����E�    �}t�}u=�=|o u4jh�`�(���u�|o   ��������2���0�E�   �E�E̋M̃��M̃}���   �U����_�$�x_�loQ�>�����E�}t�UR�0�����lo�~�poP�z>�����E�}t�MQ��/�����po�T�toR�O>�����E�}t�EP�/�����to�)�xoQ�$>�����E�}t�UR�/�����xo�E������   �j �c����Ã}� t��   ��   �}t�}t�}t��   �4&���E؃}� u�   �E؁x\�BuIhZ  h�j��NQ�$�����U؉B\�E؃x\ t��NQh�B�U؋B\P�34������j�M؋Q\R�EP�H  ���E��}� u�L�M��Q�U�}t5�E��H;Mu*�U��E�B�M����M���Nk��E�P\9U�r��ˋE��   �M�MȋUȃ��Uȃ}�w�E����_�$��_����x3�t	�E�   ��E�    �EĉEЃ}� u!h��j h�  h0�j��)������u̃}� u.�hH���    j h�  h0�h�h���=������������M�d�    Y_^[��]Ð]\]�]2]�] �I �^�^     ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h*h"�d�    P���SVW�XD1E�3�P�E�d�    j �g)�����E�    �} u!�E�lo�E܋Q�:�����E��E�   ��E�po�U܋P�:�����E��E�   �}� t�}�t
�_W���M܉�E������   �j �`����Ã}� u3���}�t
�U�R�U���   �M�d�    Y_^[��]� ��������������������������������������������������������������������̋�U��j�h(*h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    �E�    �E�EċMă��Mă}���   �U����d�$��d�E�lo�MЋ�U�E؃��E��  �E�po�MЋ�U�E؃��E���   �E�to�MЋ�U�E؃��E���   �E�xo�MЋ�U�E؃��E��   �f!���E��}� u�����  �M��Q\R�EP��  �����EЋMЋ�U��   �x3�t	�E�   ��E�    �M��Mȃ}� u!h��j h�  h0�j��%������u̃}� u1�YD���    j h�  h0�h,�h���9��������6  �E�P�:8�����E�}�u3��  �}� uj�>(���}� t
j �&�����E�    �}t�}t�}u,�M��Q`�U܋E��@`    �}u�M��Qd�ŰE��@d�   �}u<��N�M��	�Uԃ��Uԡ�N�N9E�}�M�k��U��B\�D    ���
�pT���MЉ�E������   ��}� t
j �]����Ã}u�U��BdPj�U���
�MQ�U���}t�}t�}u�U��E܉B`�}u	�M��ỦQd3��M�d�    Y_^[��]�Jb�b�b�bgb�b ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M��Q;Ut�E����E���Nk�M9M�s�ً�Nk�U9U�s�E��H;Mu�E���3���]������������������������������������̋�U��toP�w5����]�����������̋�U���yU����d]�����������������̋�U���YU����`]�����������������̋�U���<�E�    �R���E��E�    �E�    �E�    �=�o ��   h���,��E؃}� u3���  h���E�P���E�}� u3��  �M�Q�&������oh���U�R��P�&������ohx��E�P��P��%������ohX��M�Q���E�U�R��%������o�=�o th<��E�P��P�%������o��o;M�tl��o;U�ta��oP��3�����Eԋ�oQ��3�����EЃ}� t8�}� t2�UԉE�}� t�U�Rj�E�Pj�M�Q�UЅ�t�U���u�E�   �}� t�E    �E�[��o;M�t��oR�3�����Ẽ}� t�ỦE�}� t,��o;E�t"��oQ�Q3�����Eȃ}� t
�U�R�UȉE衄oP�03�����Eă}� t�MQ�UR�EP�M�Q�U���3���]������������������������������������������������������������������������������������������������������������������������������������������������̋�U���<�EԉE�3Ƀ} ���MЃ}� u!hmj h�   h�j�������u̃}� u1�>���    j h�   h�hЭhm�h3��������T  3��} ���Ẽ}� u!h\lj h�   h�j�)������u̃}� u1�=���    j h�   h�hЭh\l��2���������   �U�U��E��@B   �M�U�Q�E�M��U��B����E�Pj �MQ�U�R�;>�����E��} u�E��   �E�H���U�J�E�x |!�M�� 3�%�   �EȋM����E���M�Qj �3�����EȋU�B���M�A�U�z |"�E�� 3ҁ��   �UċE����U�
��E�Pj �2�����EċE���]��������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�X.������]������������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�)%������]����������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�UR��'������]������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�&������]����������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�g$������]��������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�EP�'������]����������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR��%������]��������������������̋�U��Q�E�E��M�Q�UR��!������]����������������̋�U��Q�E�E��M�Q�UR�������]����������������̋�U��Q�E�E��M�Q�UR�EP�x������]������������̋�U��Q�E�E��M�Q�UR�EP�/������]������������̋�U��Q�E�E��M���E����E���t��E�+E������]����������������̋�U���(�} t�} v	�E�   ��E�    �E�E�}� uhx�j jh�j�v������u̃}� u0��8���    j jh�h`�hx��N.�����   �X  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9�Hs��H�U��	�E���E�M���Qh�   �U��R��C����3��} ���E��}� uhЗj jh�j�������u̃}� u0�/8���    j jh�h`�hЗ�-�����   �  �U�U��E�E��M��Uf�f��M���E����E��M���M��t�U����U�t�˃}� ��   3��Mf��}�tJ�}���tA�}v;�U��9�Hs
��H�E��	�M���M��U���Rh�   �E��P��B���������t3�t	�E�   ��E�    �E܉E�}� uhX�j jh�j�������u̃}� u-�7��� "   j jh�h`�hX��e,�����"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9�Hs��H�U���E+E����M+ȉM؋U���Rh�   �E+E��M�TAR��A����3���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � �����������������������U��WV�u�M�}�����;�v;���  ��   r�=Py tWV����;�^_u^_]������   u������r*��$��s��Ǻ   ��r����$��r�$��s��$�8s��r�rs#ъ��F�G�F���G������r���$��s�I #ъ��F���G������r���$��s�#ъ���������r���$��s�I �s�s�sxspshs`sXs�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��s���s�s�s�s�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�@u�����$��t�I �Ǻ   ��r��+��$�Dt�$�@u�Ttxt�t�F#шG��������r�����$�@u�I �F#шG�F���G������r�����$�@u��F#шG�F�G�F���G�������V�������$�@u�I �t�tuuuu$u7u�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�@u��PuXuhu|u�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��� y    ����� y3�]�������������������̋�U��E���#Py� y� y]�������������������U���������$�\$�   ��fD$f=p�f��fT���fs�,f�� fV�f��%�   ��%�  �Y<��f,���f(4����  +у�ʁ�   ���  �    �� fn�f��fs����f����fs�&f�� fT%p�%�   ��%�  �Y� ��Y,� ��fX4��fV%���X�fT���fs�f�� f���\�f=��%�  ��%�  �Y,� ��Y� �fX4�0�fT��\��X����Y��Y��Y��\��Y����\��X�fL$f���\��\�f��f���\����X��\��\�f�%�  =�  �  ���  -�?  º�@  +�-p<  Ё�   ���  �\��\�f%��fT�fT��\�fWҺ`@  f�����Y��\��\��Y��Y�f(@��Y��-��Y�f(P��X�fp���X�� +��� �-�� �� ��  ȃ��ခ��� �X����X`�fY��\`�fY��\�����f(�`�f(5��fY�fX�fp���Y�fW���?  �X�f���X�f%��fn��YT$�Y�fs�-fp�Df(=���X�fY��X�f�fY��Y�fY�fX�fY��Y�fp���Y�fp���Y��Y��XŃ��X��X��X�fD$�D$���fL$f��f~���fT�fs� f~Ɂ�  ���   ��� �  �� �  �ځ��  fs�4fVӹ�  fn�fs�f��f��f��f��fv�f�ʁ��  ���  ��  %�   =�   ��  fL$fT$��  fn�fT��fs�4f��f��f��fv�f��%�   �� ȁ�   ��r^�� fp�f���&���f|$fd$f~�fs� f~���%���=  ���  ��  �� ��  �  �    fW���C  f��f=p�f���Y�f~�fs� f~��� tRfT���fT��fs�,f�� fV�%�   ��%�  �Y<��f,���f(4���> �\����Ё������ u��T$��   ��� t1��#��  ��fn�fs� f��fT$�^ʺ   �  ��#��� ��   ���fp�fW�fT�fv�f�Ɂ��   ���   ��   f���� �  �� ��   %�   =�   uefL$fT$��  fn�fT��fs�4f��f��f��fv�f��%�   =�   t#fL$f��% �  �� t��������fL$f��% �  �� �G  ���fL$f��% �  �� �+  ����X��ĺ�  �  fT$f~�fs� f~ҁ����¹    �� �����f��f��Yɺ   �H  fd$fT$fp�fW�fT�fv�f��%�   =�   ��   f~��� u fs� f~��  �?��   ��  �u���fp�fW�fT�fv�f��%�   =�   uUf��fd$% �  ��  �у� ��   �� tf��%�  =�?  r���f��%�  =�?  s��������X��º�  �cf~�fs� f~��������f���   �� t:f~�   %���=  �w%r�� w��fD$�D$���f��   ��fD$�T$�ԃ��T$���T$���$�	���D$��Ã� ~(=   �<  V�Ѓ��� � ��   ��W��?  �&= ����  V�Ѓ����   � � W�    �X����X`����� fY��\`�fY��\�����f(�`�f(5��fY�fX�fp���Y��X��X�f%��fnʁ�� �������� �fW���?  f���YT$�Y�fs�-fp�Df(=���X�fY��X�f�fY��Y�fY�fX�fY��Y�fp���Y�fp���Y��Y�fn�fs�-fn�fv�f���X��X�fT��X�fW�fv�f���\����X�fT�f��_�\��X��XÃ� N^�Y��Y��X��Y��X�f��%�  �   =�  �����   �� ������fD$�D$���^�X��Y��Y��X�f��%�  �   =�  ������   �� �������fD$�D$���f�fn��Y�fs�-fV��   �����   �� tf���Y ��e���f ��Y��T���fp�DfY�f��%�  ��@  +�-p<  Ё�   ������=   �r �ɀ� fn�fs�-��fD$�D$���fd$f�����  ���?  f��3�% �  �� �-����K�����$    ��$    �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ƅp����
�uK�����ƅp����2������;  ������a���t��=,it�����)����@u��
�t���2  �F  �t2��t��������(  �  �����-�Lƅp����������ݽ`������a���Au����ƅp������-�L�
�uS��������
�u������  ��   ����
�u���u
�t���ƅp����-�L��u�
�t��������  ���(  X��ݽ`������a���u���-�L
�t���ƅp����W  �����-�Lƅp����
�u����-�L������-�L�ٛݽ`������a���Au�������ݽ`������a���������ݽ`�������������ٛ���u����L�����ٛ���t�   ø    ���   ��V��t��V���$���$��v�������f���t^��t�C  �����������������������������������������������������������������������������������������������������������������������������������������̀zuf��\���������?�f�?f��^���٭^����LM�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^����LM�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp����DM���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-0M��p��� ƅp���
��
�t�������������������������������������������������������������������������������������������������������������������������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�2�����E�f�}t�m���������������������������������������������������ËT$��   ��f�T$�l$é   t�   �����   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   ���Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t�W��Z���0��Z��,$Z����������������������   s��������������������������   v��������������������������������������������������������������������������������������������������������̋�U���,�E�    ���]����Au
�E���]���E�]��E��]��}  �u@�} u:���]�����z�E��W�����]�����Au	�M�����U����%  �}  ��uK�} uE���]�����z	�E����+���]�����Au�M��W���U��W��E�   ��   �}  �u@�} u:���]����z�E��W�����]����Au	�M�����U����   �}  ��u�} uy���E�$�_������E����]����z&�}�u��W���]��	��W�]܋E�E���3���]����Au �}�u�X�]�����]ԋM�E����U����E���]����������������������������������������������������������������������������������������������������������̋�U������E�$�:�����%�   t3��\���E�$�	������]��E�]�����Dz9�E�5H.���$��������E�5H.������Dz	�   ���   �3���]��������������������������������������������̋�U���X�E�E��} t�} v	�E�   ��E�    �MĉM�}� uhX�j jOh��j���������u̃}� u0�B���    j jOh��h��hX�������   �{  �E�  �}�tI�}���t@�}v:�M��9�Hs��H�U��	�E���E��M�Qh�   �U��R�(#�����}����E�uh|�j jVh��j�	�������u̃}� u0����    j jVh��h��h|��������   ��  3҃} �U�}� uhX�j jZh��j��������u̃}� u0�%���    j jZh��h��hX��{�����   �^  �M3҃y �U��}� uh$�j j^h��j�:�������u̃}� u0����    j j^h��h��h$�������   ��  �M�y |�U�z	�E�   ��E�    �E��E܃}� uh��j jch��j��������u̃}� u0�:���    j jch��h��h��������   �s  �U�z |�E�x	�E�   ��E�    �M��M؃}� uh8�j jhh��j�6�������u̃}� u0����    j jhh��h��h8�������   ��  �E�x |�M�y;	�E�   ��E�    �U��Uԃ}� uh��j jlh��j��������u̃}� u0�6���    j jlh��h��h���
�����   �o  �M�9 |�U�:;	�E�   ��E�    �E��EЃ}� uhH�j jph��j�4�������u̃}� u0����    j jph��h��hH��
�����   ��  �U�z��   �E�H�U�B��Y+�Y�U;J}]�E�H��l  ��  �yI���A��u�U�Bl  ��d   ����u�U�Bl  ���  ����u�U�zu�E�x	�E�   ��E�    �M��M̃}� u!hp�j h�   h��j�5�������u̃}� u3����    j h�   h��h��hp��
	�����   ��  �E�x |�M�y	�E�   ��E�    �U��Uȃ}� u!h��j h�   h��j��������u̃}� u3�/���    j h�   h��h��h��������   �e  �M�Qk��U��E�Hk��M��E�    ��U���U�E����E��}�}%�M�M�U������M�M�U���4��B�ËM�� �U����U��E��  �M����M��U�BP�M�Q�  ���E��U�� �E����E��M�QR�E�P�  ���E��M��:�U����U��E�HQ�U�R�Z  ���E��E�� :�M����M��U�P�M�Q�6  ���E��U�� �E����E��M�A��d   ����P�U�R�  ���E��E�@��d   ��R�U�R��  ���E��E�� 
�M����M��U�� 3���]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E��
   ����0�U��E���E�E��
   ����0�E��M���M�E]������������������������������̋�U����E��o�E�    ������E�}� t9�E�x< u'h�   h��jjj�������M�A<�U�z< t	�E�H<�M��U��U��EPj�M�Q��%�����E��}� t3���E���]���������������������������������������̋�U���0VW�E�    �E�    �E�    �E�    3��} ���E��}� uhp�j jEh��j���������u̃}� u0�`���    j jEh��h��hp�������   �  j$h�   �UR�����3��} ���E܃}� uh��j jHh��j�e�������u̃}� u0�����    j jHh��h��h���=�����   �  �U�U؋E؃x |�M؃9 s����    �   ��  �U�UԋEԃx|"�Mԁ9�o@�v�m���    �   �  �����j jRh��h��hl��U�R�h�����P�[�����j jSh��h��h4��E�P�����P�3�����j jTh��h��h���M�Q������P�������U�UЋEЃx ��   �MЁ9�� ��   �E���M�1+��Au�E�M�Q�UR�|�����E�}� t�E���  �}� tO�EP�������t?�E���M�+ȋE�M�E�M�Q�UR�1�����E�}� t�E��  �E�@    �z  �MQ�UR������E�}� t�E��[  �}� t7�EP�������t'�M���ȋ�E�E��+��M�u�U�B    ��E� ��ȋ�E��+��M�u�j j<�U�R�E�P�'����M��U�: }�E���<�U�
�E��<�M�� �E�M�U�B�����j j<�E�P�M�Q�������u�}�j j<�U�R�E�P������M�A�U�z }!�E�H��<�U�J�E��<�M�� �E�M�U�B�����j j<�E�P�M�Q�������u�}�j j�U�R�E�P�]����M�A�U�z }!�E�H���U�J�E���M�� �E�M�j j�U�R�E�P�N����E�U�}� |D�}� v<�M�U�B���   ���E�P�M�UJ�E�H�M�UJ�E�H�   �}� ��   |
�}� ��   �M�Q�E�D��   ���E�P�M�UJ�E�H�M�y @�U�B���M�A�U�E�H��m  �E�P�M�A   �U�B���M�A��U�EP�M�Q3�_^��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��������E��}� u3�� �EP�M�Q�W������E��}� t3���E���]�������������������SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� ����������������������������������������U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�   ���E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�������E�}���]��������������������������������������������������U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]��������������������������U�������$�~$�   ��fD$f%pf�fW�fx��fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU�
fV�f($������X��\��Y��Y��Y����X��^�f(f-�\�fs�?��fs�?�Y�fp�Df5 �Y��Y���fW��Y�f\%��Y��X��Y��\�fp���X��\��\�fD$�D$���-�  ��A�-  fs�&fs�&f��fU��\����Y��X�fV��\��Y����\��Q�%�   ������fT�fs�f��fV�fn�fp� ����  ��Y<��
�Y��Y��Y��\�fT��X��\��X�f-�\��X�f(�^�f fXհ����Y��Y��Y΃��Y��Y��X�f���Y��X��X�% �  f����fp���X��\��X��X��X�fW�fD$�D$����;  = 8  ��   f�f(50f�f(@f(%PfY�f(-���fY�fY�fY����Y�fX�fY��Y�fX�fp��fY�fp���\�fp���\��\��\��\��\��X�fD$�D$���-�;  ����   fW�fT=pf%�f(0�Y�f(@�\�f(Pfp�D�Q�fY�fp�Df��fY�fX�f�fY�����Y�fX�fp�D�Y�fT�fY�fT�fp�D�\��X��Y��\��\��Y�fp���\��^��fX�fY�fp���X�% �  f��fp���X��X��X��X�fW�fD$�D$����� = � ��   f~�fs� f~�������  �?+���� ��   fT$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��:   ��fD$�T$�ԃ��T$���T$�$����fD$����fD$�D$���f������fn�fp� f�f�fT�fT��X�fD$�D$���f�f��X�fD$�D$���fW��Xƺ�  �J��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�b�������tj�S�������u#�=Hiuh�   �c����h�   �V����]�������������������������̋�U����E�    �	�E����E��}�s�M��U;�pMu��ރ}��Q  �}�   t0�}�   t'�}t!�E���tMQj j j j���������u�j��������tj��������uT�=HiuKj����E�}� t5�}��t/j �U�R�E���tMQ�����P�U���tMP�M�Q���  �}�   ��  �E��o�U���o�  +E�M�M�j h�   h�#h�#h�"h�"h  h�o������P�"������U�Ƃ   h  �E�Pj �0���u4j h�   h�#h�#h "h�!�M�Q�U�R�@�����P��������E�P����������<vT�M�Q������U��DŉE�j h�   h�#h�#hP!jhH!�M�+M�U�+�R�E�P�n�����P�g�����j h�   h�#h�#h� ht-h  h�o�������P�1�����j h�   h�#h�#h��M���tMRh  h�o������P�������h  h�h�o�k������]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�    �	�E����E��}�s�M��U;�pMu�E���tM���3���]�������������������������������̋�U���   �XD3ŉE�}��  �E�E���p����M�ǅd���    ǅh����   j ��h���R�E�P�MQ�UR�EP��������l�����l��� ��   �����zt�  j j j �MQ�UR�EP���������h�����h��� u��   j\h@%jj��h���Q�s������E��}� u��   ǅd���   j ��h���R�E�P�MQ�UR�EP�v�������l�����l��� u�   jgh@%jj��l���Q�������U���E��8 u�]j jjh�$h�$h$��l�����Q�U�R��l���P�M��R�P�����P�I�������d��� tj�E�P������3���   ��d��� tj�M�Q������������   ��   �} ��   ǅT���   �U��\���j ��T���Phts�MQ�UR�EP���������u����   ��\���� ǅ`���    ���`�������`�����`���}L��`����Ets��[�����[���R�6�������t!��\����k�
��[����DЋ�\�������3������M�3��������]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�|s]�����������������̋�U��j�hH*h"�d�    P���SVW�XD1E�3�P�E�d�    �E������E�    j�0�������u����E  j�������E�    �E�    �	�E���E�}�@��  �M�<� x �%  �U�� x�E��	�M؃�@�M؋U�� x   9E���   �M��Q����   �E؃x ucj
��������E�   �M؃y u0h�  �U؃�R���������u	�E�   ��E؋H���U؉J�E�    �   �j
������Ã}� u+�E؃�P�p��M��Q��t�E؃�P�t��2����}� u-�M��A�U�������E����M�U�+� x��E��������}��t��   ��   h�   h|%jj@j � ������E؃}� ��   �E�M؉� x��w�� ��w�	�E؃�@�E؋M�� x��   9U�s#�E��@ �M�������U��B
�E��@    뿋M����M܋U����E܃����� x�D�U�R��������u�E������������E������   �j�o����ËE܋M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�} ��   �E;�w��   �M���U������ x�<�um�=HiuB�M�M��}� t�}�t�}�t�(�URj��4���EPj��4���MQj��4��U���E������ x�U�3����$���� 	   �"����     �����]�����������������������������������������������������������̋�U��Q�} ��   �E;�w��   �M���U������ x�L����   �U���E������ x�<�th�=Hiu<�U�U��}� t�}�t�}�t�"j j��4��j j��4��
j j��4��E���M������ x�����3�������� 	   �����     �����]������������������������������������������������������������̋�U����}�u�����     ����� 	   ����2  �} |�E;�ws	�E�   ��E�    �M�M��}� u!h�fj h:  h�%j��������u̃}� u<�5����     �!���� 	   j h:  h�%h�%h�f�t���������   �E���M������ x�D
������؉E�u!h<fj h;  h�%j��������u̃}� u9�����     ����� 	   j h;  h�%h�%h<f������������U���E������ x���]����������������������������������������������������������������������������������������������̋�U��j�hx*h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    �E� �E��t
�M�� �M�U�� @  t�E��   �E�M��   t
�U���U�EP����E��}� u���P����������q  �}�u�M��@�M���}�u
�U���U������E؃}��u�����    �����     ����#  �E�    �EP�M�Q�l������U���U�E����M؃����� x�E�D
�M����U؃����� x�L$�ဋU����E؃����� x�L$�E����M؃����� x�D
$$�M����U؃����� x�D$�E�   �E������   �K�}� u8�U����E؃����� x�T����E����M؃����� x�T�M�Q�������Ã}� t�U؉U���E������EԋM�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h�*h"�d�    P���SVW�XD1E�3�P�E�d�    �E���M����� x�M��E�   �U��z uaj
�~������E�    �E��x u.h�  �M���Q��������u�E�    �U��B���M��A�E������   �j
�K����Ã}� t!�U���E������ x�TR�p��E�M�d�    Y_^[��]������������������������������������������������������������������������̋�U��E���M������ x�D
P�t�]������������������������̋�U��j�h�*h"�d�    P�ĄSVW�XD1E�3�P�E�d�    �e��E�    �E�P�<��E������,�   Ëe�ǅ|��������E�������|����  �E�����h�   hX&jj@j �������E��}� u�����  �M�� x��w    �	�U���@�U�� x   9E�s^�M��A �U�������E��@
�M��A    �U��B$$��M��A$�U��B$$�M��A$�U��B%
�E��@&
�M��A8    �U��B4 ��E҅���  �}� ��  �Mԋ�U��Eԃ��E��M�M��M��}�   }�U���x����
ǅx���   ��x����E��E�   �	�M����M���w;U���   h�   hX&jj@j �������E��}� u��w�E��   �M��U��� x��w�� ��w�	�M���@�M��U��� x   9E�sP�M��A �U�������E��@
�M��A    �U��B$$��M��A$�U��B%
�E��@&
�M��A8    �U��B4 ��,����E�    ��E����E��M����M��U����U��E�;E���   �M��9���   �U��:���   �E����tx�U����u�M��R�����t]�E����M������ x�M��U��E���
�U��E���Jh�  �U���R�u�������u����k  �E��H���U��J�9����E�    �	�E����E��}��,  �M��� x�M��U��:�t�E��8���   �M��A��}� uǅt���������U�����҃����t�����t���P���E��}����   �}� ��   �M�Q����E��}� tt�U��E���M����   ��u�U��B��@�M��A��U����   ��u�E��H���U��Jh�  �E���P�Y�������u����R�M��Q���E��P��M��Q��@�E��P�M��������U��B�   �M��A�������wR�8�3��M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �	�E����E��}�@}y�M��<� x tg�U��� x�E��	�M���@�M��U��� x   9E�s�M��y t�U���R�l���j�E��� xQ�V������U��� x    �x�����]���������������������������������������������������̋�U���@SVW�E�    �E�    �E�    �E-l  ��F|�M��l  ��L  ~������    �������  �U��l  �U�}|�}~�����    ��������  �} |�}~�~����    �������  �} |�};~�\����    �������  �} |�};~�:����    �������{  �}|[�E�M��Y+�Y;U}X�E%  �yH���@��u�E��d   ����u�El  ���  ����u�}u�}~������    �������  �U�E�Y�E��M��  �yI���A��u�E��d   ����u�El  ���  ����u�}~	�U����U��E���F�� j hm  RP�����ȋ�E���������E����d   ��+��E+  ���  ���D���E���j jVQ�����ȋ�E���M��u�j j<�U�R�E�P�����ȋ�E���j j<VQ�y����ȋ�E���M��u��I���j h�   h�&h�&hl��U�R������P������j h�   h�&h�&h4��E�P�������P�w�����j h�   h�&h�&h���M�Q�������P�L������E��E��M�ʉE��MċU��U�E�E��M���M܋U�UԋE�EЋM�M̃} t�} �u(�}� t"�U�R���������t�E��E��M�ʉE��MċE��U�_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h�*h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    �E������E�    3��} ���EЃ}� uh�'j jhhH'j��������u̃}� u.�?����    j jhhH'h8'h�'�����������   �U�UԋEԃ��EԋMԋQ��U��E�    �E�    j �E�Pj@�MQ�UR�E�P�M�Q��  ���E��E������   �Q�}� tJ�}� t8�U����E؃����� x�T����E����M؃����� x�T�M�Q�?�����Ã}� t�c����U�������E؋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������̋�U��j�h�*h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    3��} ���E܃}� u!hl(j h�   hH'j���������u̃}� u3�j����    j h�   hH'hH(hl(�������   �  �U�����3��} ���E؃}� u!h�'j h�   hH'j�s�������u̃}� u3������    j h�   hH'hH(h�'�H������   �  �} to�U�������҃��U�u!h�'j h�   hH'j���������u̃}� u3�����    j h�   hH'hH(h�'��������   �   �E�    �MQ�UR�EP�MQ�UR�EP�M�Q�)  ���E��E������   �[�}� tT�}� t@�U����M������� x�L����U����U������� x�L�M�R茻����Ã}� t	�E� �����E�M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���   �E�    �E� �E�    �E�   �E�    �E%�   t�E�    �E���E�   �E� j h�   hH'h�*h�*�M�Q�������P�������U�� �  u/�E% @ t�M��ɀ   �M���}� �  t�U��ʀ   �U��E���E�t�}�t�}�t6�@�E�   ���   �M��t�U��   t	�E�   ���E�   @�   �E�   ��   ������     �E� ����3�t	�E�   ��E�    �U��U��}� u!h@*j h  hH'j��������u̃}� u3�����    j h  hH'h�*h@*��������   �  �M�M��U����U��}�pw_�E�����$����E�    ��   �E�   ��   �E�   �   �E�   �   �}�   �u	�E�   ��E�    �   ������     �U�����3�t	�E�   ��E�    �M��M��}� u!h�)j h2  hH'j��������u̃}� u3�����    j h2  hH'h�*h�)��������   �  �E%   �E��}�   7�}�   tK�}�   �}�   t]�}� t3�}�   t6�d�}�   tO�Y�}�   t,�}�   t/�}�   t�<�E�   �   �E�   �   �E�   �   �E�   �   �E�   �   ������     �M�����3�t	�E�   ��E�    �E��E��}� u!h@*j hT  hH'j��������u̃}� u3�b����    j hT  hH'h�*h@*�������   �  �E�   �U��   t�(o��#E%�   u�E�   �M��@t �U��   �U�E�   �E��M���M�U��   t�E�   �E�M�� t�U��   �U���E��t�M��   �M��|����U��E�8�u+�����     �M������w����    �l���� �
  �U�   j �E�P�M�Q�U�R�E�P�M�Q�UR�@��E��}���  �E�%   �=   ���   �M����   �U�������U�j �E�P�M�Q�U�R�E�P�M�Q�UR�@��E��}��u^�E����U������� x�T����E����E� ������ x�T���P�F�����������U���	  �^�E����U������� x�T����E����E� ������ x�T���P�������'�����U��g	  �E�P����E�}� ��   �E�    �M����E������� x�D
����M����M�	������ x�D
����E��E�P�d������M�Q����}� u�����    ������U���  �}�u�E���@�E���}�u
�M����M��U�R�E�Q��������U����U��E����U������� x�U��T�E����U������� x�T$�​E����E� ������ x�T$�U���H��   �E�%�   ��   �M����   jj��U�P��������Eă}��u/製���8�   t�M�R����������� �E��  �   �E� j�M�Q�U�P�-�������u?�Mσ�u6�EęRP�U�P�#��������u�M�R�P���������� �E��_  j j �M�R�.������Eă}��u�E�Q�������������U��'  �E�%�   �;  �M�� @ u'�Uȁ� @ u�E @  �E��Mȁ� @ M�M�U�� @ u!h`)j h,  hH'j��������u̋M�� @ ��|�����|���   2��|���   ti��|��� @  t@��|���   t:��|��� @ t.�M��|��� @ t7��|���   t1��|��� @ t%�'�E� �!�U��  ��  u�E��
�E���E��E%   �5  �E�    �E�    �E�    �M���@��  �U���   ���x�����x���   @t-��x���   �t��x���   ���   �  �E�   �  �EЉ�t�����t�������t�����t�����   ��t����$���jj j �E�Q��������l�����p�����l����p���tPj j j �E�Q�d�������d�����h�����d���#�h������u�E�Q�������������U���  ��E�   ��   �EЉ�`�����`�������`�����`�����   ��`����$���jj j �E�Q���������X�����\�����X����\���tWj j j �E�Q��������P�����T�����P���#�T������u�E�Q�/������������U��>  �E�   ��E�   ��E�   �}� ��  j�E�P�M�R�������E��}� ~2�}�u,3�u!h,)j h�  hH'j���������u��E�    �U���L�����L����t��L���t=��L���t"��   �E�Q�w������F�����U��  �}�﻿ u	�E���   �E�%��  =��  uJ�M�R�9�����3�u!h�(j h�  hH'j�[�������u�������    �E�   �  �U�����  ����  u>j j�E�Q��������Eă}��u�U�P�������������M���  �E��8j j �U�P�������Eă}��u�M�R�������T���� �E��  �}� ��   �E�    �E�    �E�    �MH�����H���t��H���t��E���  �E�   ��E�﻿ �E�   �U�;U�~U�E�    �E�+E�P�M��T�R�E�Q��������E��}��u�U�P�������������M���  �U�U��U�룋E����U������� x�U���D$$�
M����M�	������ x�D
$�E%   ����؋M����M�	������ x$���L
$��
ȋU����U������� x�L$�M���HuH�U��t@�E����U������� x�T�� �E����E� ������ x�T�U���   ���   ���   �E����   �M�Q����U�������U��E�   j �E�P�M�Q�U�R�E�P�M�Q�UR�@��E��}��uk���P�������E����U������� x�T����E����E� ������ x�T�U�P�������������M��"� �U����M������� x�M���E���]Ë�_�k�w������� �I ����u�u�������1�1��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E������E�E��M����M��U��B��E��E�    j �M�Q�U�R�EP�MQ�UR��������E�}� t	�E�������E��E�E��]������������������������������̋�U��j�EP�MQ�UR�EP�MQ������]�����������̋�U��j�h+h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    �E������E�    3��} ���EЃ}� uh�'j jhhH'j�-�������u̃}� u.�����    j jhhH'h�*h�'�����������   �U�UԋEԃ��EԋMԋQ��U��E�    �E�    j �E�Pj@�MQ�UR�E�P�M�Q��  ���E��E������   �Q�}� tJ�}� t8�U����E؃����� x�T����E����M؃����� x�T�M�Q诤����Ã}� t������U�������E؋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������̋�U��j�h8+h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    3��} ���E܃}� u!hl(j h�   hH'j�X�������u̃}� u3������    j h�   hH'h�*hl(�-������   �  �U�����3��} ���E؃}� u!h�'j h�   hH'j��������u̃}� u3�e����    j h�   hH'h�*h�'踺�����   �  �} to�U�������҃��U�u!h�'j h�   hH'j�n�������u̃}� u3������    j h�   hH'h�*h�'�C������   �   �E�    �MQ�UR�EP�MQ�UR�EP�M�Q�)  ���E��E������   �[�}� tT�}� t@�U����M������� x�L����U����U������� x�L�M�R�������Ã}� t	�E� �����E�M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���   �E�    �E� �E�    �E�   �E�    �E%�   t�E�    �E���E�   �E� j h�   hH'h�*h�*�M�Q�h�����P�$������U�� �  u/�E% @ t�M��ɀ   �M���}� �  t�U��ʀ   �U��E���E�t�}�t�}�t6�@�E�   ���   �M��t�U��   t	�E�   ���E�   @�   �E�   ��   �j����     �E� ����3�t	�E�   ��E�    �U��U��}� u!h@*j h  hH'j脣������u̃}� u3�����    j h  hH'h�*h@*�Y������   �  �M�M��U����U��}�pw_�E������$����E�    ��   �E�   ��   �E�   �   �E�   �   �}�   �u	�E�   ��E�    �   �h����     �U�����3�t	�E�   ��E�    �M��M��}� u!h�)j h2  hH'j肢������u̃}� u3�����    j h2  hH'h�*h�)�W������   �  �E%   �E��}�   7�}�   tK�}�   �}�   t]�}� t3�}�   t6�d�}�   tO�Y�}�   t,�}�   t/�}�   t�<�E�   �   �E�   �   �E�   �   �E�   �   �E�   �   �6����     �M�����3�t	�E�   ��E�    �E��E��}� u!h@*j hT  hH'j�P�������u̃}� u3�ҿ���    j hT  hH'h�*h@*�%������   �  �E�   �U��   t�(o��#E%�   u�E�   �M��@t �U��   �U�E�   �E��M���M�U��   t�E�   �E�M�� t�U��   �U���E��t�M��   �M�������U��E�8�u+�����     �M����������    �ܾ��� �
  �U�   j �E�P�M�Q�U�R�E�P�M�Q�UR�D��E��}���  �E�%   �=   ���   �M����   �U�������U�j �E�P�M�Q�U�R�E�P�M�Q�UR�D��E��}��u^�E����U������� x�T����E����E� ������ x�T���P趝�����������U���	  �^�E����U������� x�T����E����E� ������ x�T���P�V�����藽����U��f	  �E�P����E�}� ��   �E�    �M����E������� x�D
����M����M�	������ x�D
����E��E�P�Ԝ�����M�Q����}� u�����    �������U���  �}�u�E���@�E���}�u
�M����M��U�R�E�Q�A������U����U��E����U������� x�U��T�E����U������� x�T$�​E����E� ������ x�T$�U���H��   �E�%�   ��   �M����   jj��U�P�C������Eă}��u/�����8�   t�M�R� ���������� �E��  �   3�f�M�j�U�R�E�Q��������u?�Ũ�u6�EęRP�E�Q���������u�U�P������荻����M��\  j j �U�P�������Eă}��u�M�R�������U���� �E��$  �M���   �8  �U�� @ u'�E�% @ u�M�� @  �M��Uȁ� @ U�U�E% @ u!h`)j h,  hH'j�Q�������u̋U�� @ ��|�����|���   2��|���   tg��|��� @  t@��|���   t:��|��� @ t.�K��|��� @ t5��|���   t/��|��� @ t#�%�E� ��E%  =  u�E��
�E���E��M��   �4  �E�    �E�    �E�    �U���@��  �E�%   ���x�����x���   @t-��x���   �t��x���   ���   �  �E�   �  �MЉ�t�����t�������t�����t�����   ��t����$��jj j �M�R��������l�����p�����l����p���tPj j j �M�R���������d�����h�����d���#�h������u�M�R�[������*���� �E���  ��E�   ��   �MЉ�`�����`�������`�����`�����   ��`����$�$�jj j �M�R�F�������X�����\�����X����\���tWj j j �M�R��������P�����T�����P���#�T������u�M�R�������n���� �E��=  �E�   ��E�   ��E�   �}� ��  j�M�Q�U�P�������E��}� ~2�}�u,3�u!h,)j h�  hH'j�l�������u��E�    �E���L�����L����t��L���t=��L���t"��   �M�R�������趷��� �E��  �}�﻿ u	�E���   �M�����  ����  uJ�U�P������3�u!h�(j h�  hH'j�ɘ������u��Q����    �E�   �  �E�%��  =��  u>j j�M�R�I������Eă}��u�E�Q�3�����������U���  �E��8j j �E�Q�������Eă}��u�U�P��������Ķ����M��  �}� ��   �E�    �E�    �E�    �UH�����H���t��H���t��E���  �E�   ��E�﻿ �E�   �E�;E�~U�E�    �M�+M�Q�U��D�P�M�R�d������E��}��u�E�Q�I�����������U���  �E�E��E�룋M����E������� x�E�$�L
$��
ȋU����U������� x�L$�M��   ����ًU����U������� x�����T$��
ыE����E� ������ x�T$�U���HuH�E��t@�M����E������� x�D
�� �M����M�	������ x�D
�E�%   �=   ���   �M����   �U�R����E�%����E��E�   j �M�Q�U�R�E�P�M�Q�U�R�EP�D��E��}��uk���P�]������M����E������� x�D
����M����M�	������ x�D
�E�Q�}������P�����U��"� �E����U������� x�U���E���]ÍI �������=� �I ��������O�O�����O������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E������E�E��M����M��U��B��E��E�    j �M�Q�U�R�EP�MQ�UR�(������E�}� t	�E�������E��E�E��]������������������������������̋�U��j�EP�MQ�UR�EP�MQ�������]�����������̋�U��} u��s    ��EP�
�������w��s   ]����������������������������̋�U���`�XD3ŉE��E� �E� �E� �E� �E� �E� �E���E��E���E���E���E���E���E���E���E��E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E���E���E���E���E���E���E���E���E���E���E� �E� �E� �E� �E� �E� �E� �E׀�=�s t��wP聡�����E���E���M��M؋U�U��}��  4�}��  ��  �E����E��}��   ��  �M�����$�l�E�-�  �E��}���  �M��$�T�E�   �E��+�U��]��E� �]��M��]ȍU�R�U؃���u軬��� "   �E�E���c  �E�   �E��+�M��]��U��]��E� �]ȍM�Q�U؃���u�o���� !   �U�E���  �E�   �E��+�E� �]��M��]��U��]ȍE�P�U؃���u�#���� "   �M�E����  �E�   �E��+�U��]��E� �]��M��]ȍU�R�U؃���u�׫��� !   �E�E���  �E�   �E��+�M��]��U��]��E� �]ȍM�Q�U؃���u苫��� "   �U�E���3  �E�   �E��+�E� �]��M��]��U��]ȍE�P�U؃��M�E����  �E�   �E��+�U�����  �E�   �E��+�E� �]��M��]��U��]ȍE�P�U؃���u����� "   �M�E���  �E�   �E��+�U��]��E� �]��M��]ȍU�R�U؃��E�E���S  �E�   �E��+�M��]��U��]��E� �]ȍM�Q�U؃���u�_���� "   �U�E���  �E�   �E��+�E� �]��M��]��U��]ȍE�P�U؃���u����� !   �M�E���  �E�   �E��+�U��]��E� �]��M��X.�U��E� �]��M��]��U��]ȍE�P�U؃���u觩��� !   �M�E���O  �E�   �E��+�U��]��E� �]��M��]ȍU�R�U؃���u�[���� !   �E�E���  �E�   �E��+�M��]��U��]��E� �]ȍM�Q�U؃���u����� !   �U�E���  �E�   �E��+�E� �]��M��]��U��]ȍE�P�U؃���u�è��� "   �M�E���k  �E�   �E��+�U��X.�E��M��]��U��]��E� �]ȍM�Q�U؃���u�g���� !   �U�E���  �E�   �E��+�E� �X.�M��U��]��E� �]��M��]ȍU�R�U؃���u����� !   �E�E���  �E�   �E��+�M��X.�U��E� �]��M��]��U��]ȍE�P�U؃���u诧��� !   �M�E���W  �E�   �E��+�U��X.�E��M��]��U��]��E� �]ȍM�Q�U؃���u�S���� !   �U�E����  �E�   �E��+�E� �X.�M��U��]��E� �]��M��]ȍU�R�U؃���u������ !   �E�E���  �E�   �E��+�M��X.�U��E� �]��M��]��U��]ȍE�P�U؃���u蛦��� !   �M�E���C  �E�   �E��+�U��]��E� �]��M��]ȍU�R�U؃���u�O���� !   �E�E����  �E�   �E��+�M��X.�U��E� �]��M��]��U��]ȍE�P�U؃���u����� !   �M�E���  �E�   �E��+�U��]��E� �]��M��]ȍU�R�U؃���u觥��� !   �E�E���O  �E�   �E��+�M��]��U��]��E� �]ȍM�Q�U؃���u�[���� !   �U�E���  �E�   �E��+�E� �M�M��U��]��E� �]��M��]ȍU�R�U؃���u����� !   �E�E���   �E�   �E��+�M��M�U��E� �]��M��]��U��]ȍE�P�U؃���u詤��� !   �M�E���T�E�   �E��+�U��M�E��M��]��U��]��E� �]ȍM�Q�U؃���u�S���� !   �U�E���M�3��'�����]Ë�����E�����)�����f�	�U���Y����\ 	
�I M��� a � e�Y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���h��  ��NP�l������E��M���  ���  ��   ���E�$蠮�����E�}� ~C�}�~�}�t�5h��  �U�R�������E��   �E�P���E�$j�������   �M�Q�E�X.���$���E�$jj�������{���E�$�b������]��E�]�����Dzh��  �U�R蚱�����E��D�B�E��� th��  �M�Q�z������E��$�"�U�R���E��$���E�$jj�o������]���������������������������������������������������������������������������������������U�������$�~$�   ��fD$f��f%�f-00f=��B  f04�Y�f84�-��X�fP4�\�f(@4�Y�fɁ�v ����?f(- 4��+���fY��\��YX4�\�fxf����\�fY�f\�f(5 4�Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-4�Y fX5�3fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���+f��f%�f����f�4�\�fL$�D$����&U���I ��������������������������������������������������������������������������������������������������������������������U�������$�~$�   ��fD$f��f%�f-00f=��B  f�>�Y�f�>�-��X�f�>�\�f(�>�Y�fɁ� v ����?f(-�>�`6���fY��\��Y�>�\�fxf����\�fY�f\�f(5p>�Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-�>�Y fX5`>fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���I��f��f=�u�Y�>fD$�D$���f�>�Y��\��Y�>fD$�D$����hT��������������������������������������������������������������������������������������������������������������������������̋�U����=$y u詟���E�    �<i�E��}� u����e  �M����t,�E����=t	�U����U��E�P�*������M��T�U���juh�Ajj�E���P�n������E�M�8o�=8o u�����   �<i�U��	�E�E��E��M������   �E�P蹧�������E��M����=��   j~h�Ajj�E�P��������M��U�: uj�8oP�5������8o    ����rj h�   hAh�@h�@�M�Q�U�R�E�Q蒚����P�!������U���U��B���j�<iP�Ӈ�����<i    �M��    �y   3���]��������������������������������������������������������������������������������������������������������������������̋�U����E�    �=$y u蒝����t h  h�sj �0�h�s�2������=�� t������t����U���E�s�E�E�M�Q�U�Rj j �E�P��   ���}����?s�}��r����w�M��U���;E�s����dh�   h�Aj�M��U���P�r�����E��}� u����8�M�Q�U�R�E��M���R�E�P�M�Q�   ���U����,o�E��0o3���]�������������������������������������������������������������������������̋�U��E�Ho]�����������������̋�U����E�     �M�   �U�U��} t�E�M��U���U�E�    �E����"u3҃}� �U��E���M�U����U��w�E����U�
�} t�E�M����E���E�M���U�E����E��M�Q�\�������t/�U����M��} t�U�E���
�U���U�E����E��M��t �}� �M����U�� t�E��	�7����M��u�U����U���} t�E�@� �E�    �M����t!�E���� t�U����	u�M����M��ߋU����u��  �} t�M�U��E���E�M����E��E�   �E�    �M����\u�E����E��M���M���U����"uH�E�3ҹ   ���u0�}� t�U��B��"u�M����M���E�    3҃}� �U��E���E�M�U���U��t$�} t�E� \�M���M�U����M��̋U����t�}� u�M���� t�E����	u�   �}� ��   �} tQ�U��P�~�������t)�M�U����M���M�U����U��E����U�
�E�M����E���E�)�M��R�-�������t�E����E��M����E��M����E��M����M��|����} t�U� �E���E�M����E�������} t�M�    �U���U�E����U�
��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�    �=�t u0�T��E��}� t��t   ������xu
��t   �=�t��   �}� u�T��E��}� u3��  �E��E�M����t�E���E�M����u	�E���E��؋M�+M������M�j j j j �U�R�E�Pj j �ؒ�E��}� tjahBj�M�Q��l�����E�}� u�U�R�P�3��	  j j �E�P�M�Q�U�R�E�Pj j �ؒ��uj�M�Q�F������E�    �U�R�P��E���   �=�tt�=�t ��   �}� u�L��E�}� u3��   �E�E��M����t�E����E��M����u	�E����E��؋M�+M���M�h�   hBj�U�R��k�����E��}� u�E�P�H�3��%�M�Q�U�R�E�P�i{�����M�Q�H��E��3���]���������������������������������������������������������������������������������������������������������������������������������������������̋�V�0���=��s���t�Ѓ�����r�^����������̋�V�����=��s���t�Ѓ�����r�^����������̋�U��Q�E�    �   ��]����������̋�U��j h   3��} ��P�\���t�=�t u3��D�����w�=�wu,h�  �O�������u��tQ�X���t    3���   ]��������������������������������������������̋�U����=�wuo�|w�E��E�    �	�M����M��U�;xw}5h �  j �E��HQ�d��U��BPj ��tQ�`��U����U�뷡|wPj ��tQ�`���tR�X���t    ��]�����������������������������������������������������̋�U��=�t u!h�Bj h(  h@Bj�5o������u̡�t]��������������������������̋�U����E�    �E�    �=XDN�@�t�XD%  ��t�XD�щ\D�   �U�R����E��E�M�3M��M��p�3E�E��Ē3E�E��l�3E�E�U�R�h��E�3E�E�M�3M�M�}�N�@�u	�E�O�@���U��  ��u�E���E�E�M�XD�U��҉\D��]���������������������������������������������������������������������̋�U��]���������̋�U��}csm�u�EP�MQ芅������3�]����������̋�U����h���E��}� u3��  �E��H\Q�UR�  ���E��}� u	�E�    �	�E��H�M�}� u3��j  �}�u�U��B    �   �P  �}�u����B  �E��H`�M�U��E�B`�M��y�   ��N�U��	�E����E���N�N9M�}�U�k��E��H\�D    �ЋU��Bd�E�M��9�  �u�U��Bd�   �   �E��8�  �u�M��Ad�   �q�U��:�  �u�E��@d�   �Z�M��9�  �u�U��Bd�   �C�E��8�  �u�M��Ad�   �,�U��:�  �u�E��@d�   ��M��9�  �u
�U��Bd�   �E��HdQj�U���U��E�Bd��M��A    �U��BP�U���M��U�Q`�����]��������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M��;Ut�E����E���Nk�M9M�s�ڋ�Nk�U9U�s
�E��;Mt3���E���]�������������������������U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP��   ���E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�wg�����E��u�}�M�����ʃ��E�]��u��}��]��������������������������������������������������������������U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�����������������������������������������̋�U����} uhpDj jdh�Cj�i������u̋M�M��U�R菜�����E��E��H��   u$�m���� 	   �U��B�� �M��A����G  �-�U��B��@t"�>���� "   �M��Q�� �E��P����  �M��Q��tH�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J�����  �E��H���U��J�E��H���U��J�E��@    �E�    �M��M�U��B%  u6������ 9E�t�������@9E�u�M�Q�^}������u�U�R�q������E��H��  ��   �U��E��
+Hy!h`Cj h�   h�Cj�g������u̋E��M��+Q�U��E��H���U��
�E��H���U��J�}� ~�E�P�M��QR�E�P��������E��q�}��t!�}��t�M����U������ x�U���E�PN�E��H�� t7jj j �U�R��������E�U�E�#E���u�M��Q�� �E��P����O�M��Q�E���E�   �M�Q�UR�E�P�`������E�M�;M�t�U��B�� �M��A�����E%�   ��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  �XD3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M��po���E�    3Ƀ} �������������� u!h�nj h  h�Ej�/e������u̃����� uF讃���    j h  h�Eh�Eh�n�y����ǅ(��������M��J�����(�����  �E�������������Q��@��   ������P�O������������������t-�������t$������������������� x������
ǅ���PN������H$�����х�uV�������t-�������t$������������������� x������
ǅ���PN������B$�� ���ȅ�tǅ���    �
ǅ���   ����������������� u!hpmj h  h�Ej�c������u̃����� uF�9����    j h  h�Eh�Ehpm�w����ǅ$��������M��Ղ����$����O  3Ƀ} �������������� u!hmj h  h�Ej�2c������u̃����� uF豁���    j h  h�Eh�Ehm�w����ǅ ��������M��M����� �����  ǅ����    �E�    ǅ����    �E�    �E�    �E��������������E���E���a  ������ �T  �������� |%��������x���������D��������
ǅ���    ���������������������������D���������������� ����� �����  �� ����$�5�E�    �M��\a��P������R�[c��������   ������P�MQ������R�l  ���E��������U���U����������؉�����u!h�Ej h�  h�Ej�sa������u̃����� uF�����    j h�  h�Eh�Eh�E�Eu����ǅ��������M�莀��������  ������R�EP������Q�  ����  �E�    �UԉU؋E؉E�M�M��E�    �E������E�    �  �������������������� ������������wK��������@5�$�(5�E����E��,�M����M��!�U����U���E��   �E��	�M����M��!  ��������*u(�EP��z�����E�}� }�M����M��U��ډU���E�k�
�������TЉU���  �E�    ��  ��������*u�MQ�zz�����EЃ}� }�E�������U�k�
�������LЉM��  ��������������������I������������.�  ��������h5�$�T5�E���lu�U���U�E�   �E��	�M����M���   �U���6u&�M�Q��4u�E���E�M��� �  �M��   �U���3u#�M�Q��2u�E���E�M�������M��S�U���dt7�M���it,�E���ot!�U���ut�M���xt�E���Xu�ǅ����    ������U��� �U���E�   �E��J
  ��������������������A������������7�  ���������5�$��5�U���0  u�E�   �E��M���  tUǅ����    �UR�n����f������������Ph   ������Q�U�R�~���������������� t�E�   �&�EP�Ux����f�������������������E�   �������U��]  �EP�!x������|�����|��� t��|����y u��N�U��E�P�%������E��P�M���   t&��|����B�E���|�����+����E��E�   ��E�    ��|����B�E���|�����U���  �E�%0  u�M���   �M��}��uǅ��������	�UЉ�������������t����MQ�Nw�����E��U���  te�}� u��N�E��E�   �M���p�����t�����t�������t�����t��p������t��p�������p����ɋ�p���+M����M��[�}� u	��N�U��E���x�����t�����t�������t�����t��x������t��x�������x����ɋ�x���+E��E��  �MQ�ov������l���踒������   3�tǅ����   �
ǅ����    ��������h�����h��� u!hPEj h�  h�Ej�}[������u̃�h��� uF��y���    j h�  h�Eh�EhPE�Oo����ǅ��������M��z��������  ��  �U��� t��l���f������f����l�����������E�   �  �E�   �������� �������U���@�U��������E��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}У   ~Bh�  hEj�UЁ�]  R�-T�����E��}� t�E��E��MЁ�]  �M���EУ   �U���U�E�H��P���`�����d����M��Y��P�E�P�M�Q������R�E�P�M�Q��`���R�TIP�l�����Ѓ��M���   t&�}� u �M��9Y��P�U�R�`IP�al�����Ѓ���������gu,�U���   u!�M��Y��P�E�P�\IQ�)l�����Ѓ��U����-u�M���   �M��U����U��E�P�������E��	  �M���@�M��E�
   �o�E�
   �f�E�   ǅ����   �
ǅ����'   �E�   �U���   t�E�0��������Q�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ��������P�����T����   �U���   t�EP��������P�����T����   �M��� tB�U���@t�EP��r��������P�����T�����MQ��r���������P�����T����=�U���@t�EP�r�������P�����T�����MQ�r����3҉�P�����T����E���@t@��T��� 7|	��P��� s,��P����ً�T����� �ډ�H�����L����E�   �E����P�����H�����T�����L����E�% �  u&�M���   u��H�����L����� ��H�����L����}� }	�E�   ��M�����M��}�   ~�E�   ��H����L���u�E�    �E��E��MЋUЃ��UЅ���H����L���t{�E��RP��L���Q��H���R�u����0��\����E��RP��L���P��H���Q�)s����H�����L�����\���9~��\����������\����E���\�����U����U��g����E�+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@t?�E�%   t�E�-�E�   �(�M���t�E�+�E�   ��U���t�E� �E�   �E�+E�+E䉅D����M���u������R�EP��D���Qj �<  ��������R�EP�M�Q�U�R�q  ���E���t$�M���u������R�EP��D���Qj0��  ���}� ��   �}� ��   ǅ,���    �U���@����E܉�<�����<�����<�������<�������   ��@���f�f������������Rj��0���P��8���Q�u������,�����@�������@�����,��� u	��8��� uǅ���������&������P�MQ��8���R��0���P�t  ���Z����������Q�UR�E�P�M�Q�R  �������� |$�U���t������P�MQ��D���Rj ��  ���}� tj�E�P��a�����E�    �|���������������M��s��������M�3��w����]Ë�'(C(�())T)�*�(�(�(|(�(�( �I �)t*�)*�* �.�*,�/v+6.�*�/(--0�/",�/�/�2   	
���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�H��@t�U�z u�E����U�
�p�E�H���U�J�E�x |&�M��E��M���   �M��U����M���UR�EP�b�����E��}��u�M�������U����M���]���������������������������������������������������̋�U��E�M���M��~!�UR�EP�MQ�	������U�:�u���]������������������������̋�U��Q�E�H��@t�U�z u�E�M�U�
�`�E�M���M��~P�U��E��MQ�UR�E�P�������M���M�U�:�u �Uk���8*u�EP�MQj?�`�������렋�]�����������������������������������̋�U��E����U�
�E��A�]��������������������̋�U��E����U�
�E��A��Q�]�����������������̋�U��E����U�
�E�f�A�]�������������������̋�U����E�    �E�    �E�H��pt	�U��pu�E�H�U3�;����'  �E�H��st�U�B��St	�E�    ��E�   �M�M��U��st�E��St	�E�    ��E�   �M��M��}� u�}� tE�U�;U�u.�E�H��  ����ًU��  �����;�u	�E�   ��E�    �E��  �E�H��dtv�U�B��itj�M�Q��ot^�E�H��utR�U�B��xtF�M�Q��Xt:�E��dt1�M��it(�U��ot�E��ut�M��xt�U��X��   �E�H��dtE�U�B��it9�M�Q��ot-�E�H��ut!�U�B��xt�M�Q��Xt	�E�    ��E�   �E��dt6�M��it-�U��ot$�E��ut�M��xt�U��Xt	�E�    ��E�   �E�;E�t3��T�M�Q��   ����ڋE%   �����;�u�M�Q�� ����ڋE�� �����;�t3���M�3�;U����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���   �XD3ŉ�X���ǅ<���    ǅ����    ǅ����    ǅp���    ǅ����    ǅx���    ǅ����    �EP��`����xR��ǅ����    ǅ����    ǅH���    ǅ����    ǅ��������ǅ��������ǅ��������ǅ|�������ǅ��������ǅ����    3Ƀ} ����8�����8��� u!h�nj h  h�Ej��G������u̃�8��� uI�Yf���    j h  h�Eh�Oh�n�[����ǅ���������`�����f��������7  �E��4�����4����Q��@��   ��4���P��z������0�����0����t-��0����t$��0�������0�������� x��d����
ǅd���PN��d����H$�����х�uV��0����t-��0����t$��0�������0�������� x��`����
ǅ`���PN��`����B$�� ���ȅ�tǅ\���    �
ǅ\���   ��\�����,�����,��� u!hpmj h  h�Ej�bF������u̃�,��� uI��d���    j h  h�Eh�Ohpm�4Z����ǅ���������`����ze��������E6  3Ƀ} ����(�����(��� u!hmj h  h�Ej��E������u̃�(��� uI�Vd���    j h  h�Eh�Ohm�Y����ǅ ���������`�����d���� ����5  ǅT���    �E������ǅH���    ���H�������H�����H����b5  ��H���u������ u�K5  ǅ����    ǅ@���    ǅ����    ǅ\���    ǅ��������ǅ����    ǅp���    �������Uǅ��������ǅ��������ǅ|�������ǅ���������E���O�����O����E���E����1  ��T��� ��1  ��O����� |%��O�����x��O����� �����X����
ǅX���    ��X�����P�����P���k�	��@�����@�����@�����@�����  �E���%��  �������u\j
������R�EP��p������~9���������$u+��H��� uh@  j ������P�m����ǅ����   �
ǅ����    �������)  j
������Q�UR�|p���������������������E��H��� ��   ������ |#���������$u������d}ǅT���   �
ǅT���    ��T�����$�����$��� u!h�Nj hP  h�Ej��B������u̃�$��� uI�sa���    j hP  h�Eh�Oh�N��V����ǅ����������`����b����������2  ������;�����~��������P������������P�����P����������   ��@�����   3�tǅL���   �
ǅL���    ��L����� ����� ��� u!h�Nj h\  h�Ej�B������u̃� ��� uI�`���    j h\  h�Eh�Oh�N��U����ǅ����������`����$a����������1  ��@�����H�����H�����.  ��H����$�\y��H��� u	������t��H���u�������u�.  ǅ����    ��`�����@��P��O���R��B��������   ��T���P�MQ��O���R�1A  ���E���O����U���U��O�������؉����u!h�Ej h�  h�Ej��@������u̃���� uI�W_���    j h�  h�Eh�Oh�E�T����ǅ����������`�����_���������0  ��T���R�EP��O���Q�z@  ���-  ǅt���    ��t�����x�����x���������������������ǅ����    ǅp�������ǅ����    �A-  ��O�����D�����D����� ��D�����D���wi��D������y�$�|y���������������D���������������3���������������"�������   ����������������������,  ��O�����*��  ������ u�EP��Y�����������^  j
������Q�UR�7l���������������������E��H��� ��  ������ |#���������$u������d}ǅ@���   �
ǅ@���    ��@������������� u!h�Mj h�  h�Ej�>������u̃���� uI�.]���    j h�  h�Eh�Oh�M�R����ǅ����������`�����]���������.  ������;�����~��������<������������<�����<����������������������� uE��������Ǆ����   ����������O������������������������������   ������P��O���Qj��������������P�p��������؉����u!h(Mj h�  h�Ej�x=������u̃���� uI��[���    j h�  h�Eh�Oh(M�JQ����ǅ����������`����\���������[-  �M*  �+������������������������Q�W���������������� }���������������������؉������������k�
��O����DЉ�������)  ǅp���    ��)  ��O�����*��  ������ u�UR�W������p����^  j
������P�MQ�Si��������|������������U��H��� ��  ��|��� |#���������$u������d}ǅ8���   �
ǅ8���    ��8������������� u!hpLj h�  h�Ej��;������u̃���� uI�JZ���    j h�  h�Eh�OhpL�O����ǅ����������`�����Z���������+  ��|���;�����~��|�����4������������4�����4�����������|����������� uE��|�����Ǆ����   ��|�������O�����������|������������������   ������R��O���Pj��|�����������R�+m��������؉����u!h�Kj h�  h�Ej�:������u̃���� uI�Y���    j h�  h�Eh�Oh�K�fN����ǅ����������`����Y���������w*  �i'  �+��|���������������������P�T������p�����p��� }
ǅp����������p���k�
��O����DЉ�p����'  ��O�����0�����0�����I��0�����0���.�B  ��0������y�$��y�U���lu�M���M��������   �����������������������   �M���6u+�E�H��4u�U���U������ �  �������   �M���3u(�E�H��2u�U���U������%����������e�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu��������   �������ǅ@���    �*����"�������� �������������   �������%  ��O�����,�����,�����A��,�����,���7��"  ��,�����(z�$��y��������0  u������   ��������������  �_  ǅ ���    ������ u�UR�PH����f��D�����  ������ |������d}ǅ(���   �
ǅ(���    ��(��������������� u!hhKj h�  h�Ej�u7������u̃����� uI��U���    j h�  h�Eh�OhhK�GK����ǅ����������`����V���������X'  ��H��� �
  �������������� uE��������Ǆ����   ����������O������������������������������   ������R��O���Pj��������������R��h��������؉�����u!h�Jj h�  h�Ej�e6������u̃����� uI��T���    j h�  h�Eh�Oh�J�7J����ǅ����������`����}U���������H&  ��   �,��������������������������P�XF����f��D�����D���Qh   ��X���R������P��U������ ����� ��� t
ǅx���   �*  ������ u�MQ�P����f��������  ������ |������d}ǅ$���   �
ǅ$���    ��$��������������� u!hhKj h�  h�Ej� 5������u̃����� uI�S���    j h�  h�Eh�OhhK��H����ǅ����������`����8T���������%  ��H��� �
  �������������� uE��������Ǆ����   ����������O������������������������������   ������Q��O���Rj��������������Q�f��������؉�����u!h Jj h�  h�Ej�4������u̃����� uI�R���    j h�  h�Eh�Oh J��G����ǅ����������`����(S����������#  �p  �,��������������������������R�!N����f��������������X���ǅ����   ��X����������  ������ u�UR��M������������  ������ |������d}ǅ ���   �
ǅ ���    �� ��������������� u!hhKj h�  h�Ej��2������u̃����� uI�eQ���    j h�  h�Eh�OhhK�F����ǅ����������`�����Q����������"  ��H��� �
  �������������� uE��������Ǆ����   ����������O������������������������������   ������R��O���Pj��������������R�md��������؉�����u!h�Ij h�  h�Ej��1������u̃����� uI�UP���    j h�  h�Eh�Oh�I�E����ǅ����������`�����P���������!  �6  �+��������������������������P��K���������������� t�������y u#��N������������P��]�����������e��������   t/�������B��������������+���������ǅ����   �(ǅ����    �������B��������������������g  ������%0  u��������   ��������p����uǅ���������p������������������������� u�MQ��J������������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!hhKj h5  h�Ej��/������u̃����� uI�eN���    j h5  h�Eh�OhhK�C����ǅ����������`�����N����������  ��H��� �
  �������������� uE��������Ǆ����   ����������O������������������������������   ������Q��O���Rj��������������Q�ma��������؉�����u!h�Ij h9  h�Ej��.������u̃����� uI�UM���    j h9  h�Eh�Oh�I�B����ǅ����������`�����M���������  �6  �+��������������������������R��H����������������%  tx������ u��N������ǅ����   ����������������������������������t���������t���������������ɋ�����+��������������i������ u��N����������������������������������������t���������t���������������ɋ�����+������������  ������ u�UR��G������������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!hhKj h�  h�Ej��,������u̃����� uI�`K���    j h�  h�Eh�OhhK�@����ǅ����������`�����K����������  ��H��� �
  �������������� uE��������Ǆ����   ����������O������������������������������   ������R��O���Pj��������������R�h^��������؉�����u!h�Ij h�  h�Ej��+������u̃����� uI�PJ���    j h�  h�Eh�Oh�I�?����ǅ����������`�����J���������  �1  �+��������������������������P��E�����������+b������   3�tǅ���   �
ǅ���    ����������������� u!hPEj h�  h�Ej��*������u̃����� uI�oI���    j h�  h�Eh�OhPE��>����ǅ����������`����J����������  �P  �������� t������f��T���f����������T����ǅx���   �  ǅt���   ��O����� ��O�����������@��������������  ��H��� ��  ������ |������d}ǅ���   �
ǅ���    ����������������� u!hhKj h�  h�Ej�)������u̃����� uI�=H���    j h�  h�Eh�OhhK�=����ǅ����������`�����H���������  �������������� uE��������Ǆ����   ����������O������������������������������   ������Q��O���Rj��������������Q�R[��������؉�����u!h�Hj h�  h�Ej�(������u̃����� uI�:G���    j h�  h�Eh�Oh�H�<����ǅ����������`�����G���������  �  ��X���������ǅ\���   ��p��� }ǅp���   �7��p��� u��O�����guǅp���   ���p���   ~
ǅp���   ��p����   ~Zh�  hEj��p�����]  R�!���������������� t ��������������p�����]  ��\����
ǅp����   ������ u#�U���U�E�H��P��������������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!hhKj h  h�Ej�'������u̃����� uI�E���    j h  h�Eh�OhhK��:����ǅ����������`����*F����������  ��H���t!h�Hj h  h�Ej�&������u̋����������������������������������������H��P���������������`����%��P��t���P��p���Q��O���R��\���P������Q������R�TIP�8�����Ѓ���������   t/��p��� u&��`����X%��P������R�`IP�}8�����Ѓ���O�����gu5��������   u'��`����%��P������P�\IQ�<8�����Ѓ����������-u!��������   ��������������������������P�R������������  ��������@������ǅ����
   �   ǅ����
   �   ǅp���   ǅ<���   �
ǅ<���'   ǅ����   ��������   t ƅ����0��<�����Q������ǅ����   �*ǅ����   ��������   t��������   ������������% �  �#  ������ u�MQ��T������������������  ������ |������d}ǅ���   �
ǅ���    �������t�����t��� u!hhKj h�  h�Ej�$������u̃�t��� uI�B���    j h�  h�Eh�OhhK��7����ǅ����������`����C����������  ��H��� �
  �������������� uE��������Ǆ����   ����������O������������������������������   ������Q��O���Rj��������������Q�U��������؉�p���u!h�Gj h�  h�Ej��"������u̃�p��� uI�qA���    j h�  h�Eh�Oh�G��6����ǅ����������`����
B����������  �R  �1����������������l�����l���R��R������������������
  ������%   �#  ������ u�MQ�R������������������  ������ |������d}ǅ ���   �
ǅ ���    �� �����h�����h��� u!hhKj h�  h�Ej��!������u̃�h��� uI�M@���    j h�  h�Eh�OhhK�5����ǅ����������`�����@���������  ��H��� �
  �������������� uE��������Ǆ����   ����������O������������������������������   ������Q��O���Rj��������������Q�US��������؉�d���u!h@Gj h�  h�Ej� ������u̃�d��� uI�=?���    j h�  h�Eh�Oh@G�4����ǅ����������`�����?���������  �  �1����������������`�����`���R�P������������������  �������� �a  ��������@�'  ������ u�UR�:��������������������  ������ |������d}ǅ����   �
ǅ����    ��������\�����\��� u!hhKj h�  h�Ej�������u̃�\��� uI�
>���    j h�  h�Eh�OhhK�]3����ǅ����������`����>���������n  ��H��� �
  �������������� uE��������Ǆ����   ����������O������������������������������   ������R��O���Pj��������������R�Q��������؉�X���u!h Jj h�  h�Ej�{������u̃�X��� uI��<���    j h�  h�Eh�Oh J�M2����ǅ����������`����=���������^  ��  �3����������������T�����T���P�8�������������������&  ������ u!�MQ�d8���������������������  ������ |������d}ǅ����   �
ǅ����    ��������P�����P��� u!hhKj h�  h�Ej�b������u̃�P��� uI��;���    j h�  h�Eh�OhhK�41����ǅ����������`����z<���������E  ��H��� �
  �������������� uE��������Ǆ����   ����������O������������������������������   ������Q��O���Rj��������������Q��N��������؉�L���u!h Jj h�  h�Ej�R������u̃�L��� uI��:���    j h�  h�Eh�Oh J�$0����ǅ����������`����j;���������5  �  �5����������������H�����H���R�c6��������������������V  ��������@�%  ������ u�MQ�*6�������������������  ������ |������d}ǅ����   �
ǅ����    ��������D�����D��� u!hhKj h  h�Ej�+������u̃�D��� uI�9���    j h  h�Eh�OhhK��.����ǅ����������`����C:���������  ��H��� �
  �������������� uE��������Ǆ����   ����������O������������������������������   ������Q��O���Rj��������������Q�L��������؉�@���u!h Jj h  h�Ej�������u̃�@��� uI�8���    j h  h�Eh�Oh J��-����ǅ����������`����39����������	  �{  �2����������������<�����<���R�,4������������������"  ������ u�EP�4����3ɉ�������������  ������ |������d}ǅ����   �
ǅ����    ��������8�����8��� u!hhKj h/  h�Ej�������u̃�8��� uI�7���    j h/  h�Eh�OhhK��,����ǅ����������`����8����������  ��H��� �
  �������������� uE��������Ǆ����   ����������O������������������������������   ������Q��O���Rj��������������Q�J��������؉�4���u!h Jj h3  h�Ej��������u̃�4��� uI�t6���    j h3  h�Eh�Oh J��+����ǅ|���������`����7����|�����  �U  �3����������������0�����0���R�2����3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�x�����|�����������   ���������������x�����������|����������� �  u(������%   u��x�����|����� ��x�����|�����p��� }ǅp���   �%�����������������p���   ~
ǅp���   ��x����|���u
ǅ����    ��W�����������p�����p�������p�������x����|�����   �������RP��|���P��x���Q��4����0�������������RP��|���R��x���P�a2����x�����|���������9~�������<�������������������������������������K�����W���+���������������������������������   t>������ t���������0t'���������������������0��������������������u��H��� u�^  ��x��� �-  ��������@t[��������   tƅ����-ǅ����   �:��������tƅ����+ǅ����   ���������tƅ���� ǅ����   ������+�����+�������,�����������u��T���Q�UR��,���Pj �_  ����T���Q�UR������P������Q�  ����������t'��������u��T���Q�UR��,���Pj0�  �������� ��   ������ ��   ǅ���    ��������(�����������$�����$�����$�������$�������   ��(���f�f������������Qj�����R�� ���P�3�����������(�������(�������� u	�� ��� uǅT��������&��T���R�EP�� ���Q�����R�  ���Z����!��T���P�MQ������R������P�W  ����T��� |'��������t��T���R�EP��,���Qj ��  �������� tj������R�f ����ǅ����    ������@��� t��@���tǅ����    �
ǅ����   ���������������� u!h�Fj h�  h�Ej�q������u̃���� uI��0���    j h�  h�Eh�Oh�F�C&����ǅx���������`����1����x����T  �������%  ��H��� �  ǅ����    ���������������������;�������  �����������������������������������������  �������$�`z���������E�������MQ�	,�����  ���������E�������MQ��!�����_  ���������E�������MQ��+�����;  ���������E�������MQ�nA�����  ���������E�������MQ�JA������   ���������E�������MQ�U+������   ���������E�������MQ�������p�����t����   3�tǅ����   �
ǅ����    ���������������� u!h`Fj h-	  h�Ej�A������u̃���� uF��.���    j h-	  h�Eh�Oh`F�$����ǅl���������`����Y/����l����'�����������T�����h�����`����0/����h�����X���3��73����]Ë��G�H�H�IgLvL8O�PZIkIII8I~I�I �I �O�PuO�P�P ��^�PdXd�U�^Q�c�[Sd�c�X�cd�s   	
{w�w�w�wx/x�xSx�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�H��@t�U�z u�E����U�
�p�E�H���U�J�E�x |&�M��E��M���   �M��U����M���UR�EP�%�����E��}��u�M�������U����M���]���������������������������������������������������̋�U��E�M���M��~!�UR�EP�MQ�	������U�:�u���]������������������������̋�U��Q�E�H��@t�U�z u�E�M�U�
�`�E�M���M��~P�U��E��MQ�UR�E�P�������M���M�U�:�u �����8*u�EP�MQj?�`�������렋�]�����������������������������������̋�U��E����U�
�E��A��Q�]������������������U���0���S�ٽ\�����=�Z t�	����8����   [����ݕz������U���U���0���S�ٽ\����=�Z t�}	����8�����8�����Z   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���ƅq����$	���   [�À�8�����=(i uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   ��O������������O����s4��O�,ǅr���   ��O������������O����v��OVW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�/����_^�E�����U���0���S�u�u�   ���ٽ\�����8�����������[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[�������������������������������������������������������������������������������������������������������������������������������������������������������������������l$�l$�D$���   5   �   t��������N u��ËD$%�  tg=�  t`�|$�D$?  %��  �D$ �l$ �D$%�  ��t��N����N���l$�����N����N���l$��ËD$D$u��ËD$%�  u��|$�D$?  %��  �D$ �l$ �D$%�  t=�  t2�D$�s*��D$�r ��������N�|$�l$�ɛ�l$������l$��Ã�,��?�$�.O����,Ã�,�����,Ã�,�����,�����,�����,�����,��|$���<$�|$ �����l$ �Ƀ�,Ã�,��<$�|$�����l$�Ƀ�,Ã�,����|$���<$�|$ �^����l$ ��,��<$�|$�J�����,��|$�<$�:����l$��,��|$�<$�&�����,��|$�����<$�|$ �������l$ �ʃ�,Ã�,��<$���|$��������l$�ʃ�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$�����Ƀ�,��|$���<$�������l$��,��|$���<$�����Ƀ�,��|$�����<$�|$ �j������l$ �˃�,Ã�,��<$���|$�K������l$�˃�,Ã�,����|$�����<$�|$ �$������l$ ��,��<$���|$�����ʃ�,��|$���<$��������l$��,��|$���<$������ʃ�,��|$�����<$�|$ ��������l$ �̃�,Ã�,��<$���|$�������l$�̃�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�h����˃�,��|$���<$�T������l$��,��|$���<$�<����˃�,��|$�����<$�|$ �"������l$ �̓�,Ã�,��<$���|$�������l$�̓�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$������̃�,��|$���<$�������l$��,��|$���<$�����̃�,��|$�����<$�|$ �~������l$ �΃�,Ã�,��<$���|$�_������l$�΃�,Ã�,����|$�����<$�|$ �8������l$ ��,��<$���|$� ����̓�,��|$���<$�������l$��,��|$���<$������̓�,��|$�����<$�|$ ��������l$ �σ�,Ã�,��<$���|$�������l$�σ�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�|����΃�,��|$���<$�h������l$��,��|$���<$�P����΃�,Ã�,�<$�|$�;�����,Ã�,�|$�<$�(�����,�P�D$%  �=  �t3��% 8  t�D$����X� �Ƀ��<$�D$�����,$�Ƀ�X� �t$X� P�D$%  �=  �t3��% 8  t�D$�k���X� �Ƀ��<$�D$�V����,$�Ƀ�X� �t$X� P��% 8  t�D$�/���X� �Ƀ��<$�D$�����,$�Ƀ�X� P��% 8  t�D$�����X� �Ƀ��<$�D$������,$�Ƀ�X� P�D$%  �=  �t3��% 8  t�D$�����X� �Ƀ��<$�D$�����,$�Ƀ�X� �|$X� P�D$%  �=  �t3��% 8  t�D$�~���X� �Ƀ��<$�D$�i����,$�Ƀ�X� �|$X� P��% 8  t�D$�B���X� �Ƀ��<$�D$�-����,$�Ƀ�X� P��% 8  t�D$����X� �Ƀ��<$�D$������,$�Ƀ�X� P��,�<$�|$������,X�P��,�|$�<$�������,X�PSQ�D$5   �   ��  �������N �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����O�Ƀ�u�\$0�|$(���l$�-$O�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�O�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$3ҋD$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���O�|$�O�<$� �|$$�D$$   �D$(�l$(���O�<$�l$$�T�����0Z�����0Z�PSQ�D$5   �   ��  �������N �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����O�Ƀ�u�\$0�|$(���l$�-$O�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�O�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$�    �D$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���O�|$�O�<$� �|$$�D$$   �D$(�l$(���O�<$�l$$�Q�����0Z�����0Z�������@��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����} uhpDj j?h(Pj��������u̋M�M��U�R�?����P�"�������u3��  � ���� 9E�u	�E�    �� ����@9E�u	�E�   �3���   �Pi���Pi�M��Q��  t3��   �E��<��t uZj[h�Ojh   ��������M����t�U��<��t u-�E����M��A�U��E��H�
�U��B   �E��@   �/�M��U����t�A�M��U��B��M��A   �U��B   �E��H��  �U��J�   ��]����������������������������������������������������������������������������������������̋�U��Q�} t'�}t!h�Pj h�   h(Pj��������u̋M�M��} tG�U��B%   t:�M�Q�p�����U��B%�����M��A�U��B    �E��     �M��A    ��]��������������������������������������̋�U��j�hX+h"�d�    P���SVW�XD1E�3�P�E�d�    �} t�} u3��   3��} ���E��}� uh�nj jMh�Pj��������u̃}� u*����    j jMh�Ph�Ph�n�������3��L�UR�������E�    �EP�MQ�UR�EP�������E��E������   ��MQ�9�����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������̋�U���<�} t�} u3��  3��} ���E܃}� uh�nj jqh�Pj���������u̃}� u-�k���    j jqh�Ph�Rh�n�������3��A  3҃} �U؃}� uhxRj jrh�Pj��������u̃}� u-����    j jrh�Ph�RhxR�^�����3���  ���3��u;EɃ��M�uh<Rj jsh�Pj� �������u̃}� u-����    j jsh�Ph�Rh<R�������3��x  �E�E�M�M�M�U�U��E�H��  t�U�B�E���E�   �}� �5  �M�Q��  ��   �E�x ��   �M�y }I�U�z }!h`Qj h�   h�Pj�[�������u̋M�Q�� �E�P�E�+E�3��u��  �M�U�;Qs�E��E��	�M�Q�UЋEЉE�M�Q�U�R�E�Q�w������U�+U�U��E�H+M�U�J�E�M�U�
�E�E�E��T  �M�;M���   �U�B%  t �MQ�@�������t�E�+E�3��u�#  �}� t�E�3��u��E�+E���M��M̋ỦU�E�P�M�Q�UR������P������E��}��u�E�H�� �U�J�E�+E�3��u�   �E�;E�v�M�M���U��UȋEȉE�M�+M�M��U�U�U�E�;E�s�M�Q�� �E�P�E�+E�3��u�h�^�M���U��EP�M�Q�k��������u�E�+E�3��u�;�U���U�E����E��M�y ~�U�B�E���E�   �MĉM�������E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q3��} ���E��}� uh�nj j)h�Rj�>�������u̃}� u+������    j j)h�Rh�Rh�n�����������U�B��]�������������������������������̋�U��j�hx+h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    j��������E�    �E�   �	�E����E��M�;����   �U�\y�<� t|�M��\y���H��   t"�U�\y��Q��������t	�U���U�}�|=�E��\y���� R�l�j�E��\y��R�������E��\y��    �Y����E������   �j�4����ËE�M�d�    Y_^[��]����������������������������������������������������������������������������������������̋�U��j�h�+h"�d�    P���SVW�XD1E�3�P�E�d�    �}�u����� 	   ����  �} |�E;�ws	�E�   ��E�    �M؉M��}� uhTj j,h�Sj���������u̃}� u.�P���� 	   j j,h�Sh�ShT����������;  �E���M������ x�D
������؉E�uhLSj j-h�Sj�S�������u̃}� u.������ 	   j j-h�Sh�ShLS�+����������   �UR�f������E�    �E���M������ x�D
��t;�MQ�������P�t���u����E���E�    �}� u�>�L����U��9���� 	   �E�����3�uh�ej jEh�Sj�}�������u��E������   ��UR�������ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h�+h"�d�    P���SVW�XD1E�3�P�E�d�    �}�u�����     �	���� 	   ����  �} |�E;�ws	�E�   ��E�    �M؉M��}� uh�fj jDh�Tj�#�������u̃}� u9�����     ����� 	   j jDh�Th�Th�f�����������/  �E���M������ x�D
������؉E�uh<fj jEh�Tj��������u̃}� u9�(����     ����� 	   j jEh�Th�Th<f�j���������   �UR�������E�    �E���M������ x�D
��t�MQ�UR�EP�B������E��?����� 	   �����     �E�����3�uh�ej jPh�Tj���������u��E������   ��EP������ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������̋�U�츐<  �����XD3ŉE��E�    �E�    �E�    �E��E�} u3���
  3Ƀ} ���M��}� uh�hj jph�Tj��������u̃}� u9�.����     �����    j jph�Th�Uh�h�p���������
  �E���M������ x�D
$�����E��M���t	�U���uo�E��������E�uhdUj jxh�Tj��������u̃}� u9�����     �x����    j jxh�Th�UhdU������������	  �U���E������ x�T�� tjj j �EP������MQ�	�������td�U���E������ x�T��   tA����EԋEԋHl3҃y �U�E�P�M���U������ x�Q�|��E�}� ��  �}� t�U�����  �x��E��E�    �E�    �E�EЋM�+M;M�}  �U�����  �E��3҃�
�U��E���M������ x�|
8 ��   �E���M������ x�D
4P��������u!h Uj h�   h�Tj�M�������u̋U���E������ x�T4�U��EЊ�M��U���E������ x�D8    j�U�R�E�P�j��������u�  �   �M��R����������   �E�+E�M+ȃ�v'j�U�R�E�P�"��������u�O  �MЃ��M��K�U���E������ x�UЊ�T4�E���M������ x�D
8   �E����E���  �j�M�Q�U�R���������u��  �EЃ��E��4�M���t	�U���u"�E�f�f�M��U�3���
���E��MЃ��M��U�����   j j j�E�Pj�M�Qj �U�R�ؒ�Eȃ}� u�f  �[j �E�P�M�Q�U�R�E���M������ x�
P����t�M�+MM�M��U�;U�}�  �����E��	  �}� tl�E�   �E�j �E�P�M�Q�U�R�E���M������ x�
P����t!�M�;M�}�   �U���U�E����E������E��   �   �M���t	�U���u{�E�P����������U�;�u�E����E������E��R�}� tG�E�   �   f�M��U�R���������M�;�u�U����U��E���E������E���t�����  �M���U������ x�L��   �k  �E�    �U����?  ǅ����    ǅ����    �E������������+M;M�  ������������������������+�=�  sz������+U;Usl�����������������������������������
u!�M���M싕�����������������������������������������������q���j �M�Q������������+�R������Q�U���E������ x�R����t �E�E��E�������������+�9M�}������E��������  �E����C  �M������ǅ����    ������+U;U�  ������������������������+ʁ��  ��   ������+E;Esu������f�f����������������������������
u&�U���U�   ������f���������������������f������f����������������c���j �E�P������������+�Q������P�M���U������ x�Q����t �U�U��U�������������+�9E�}������E���������  �U������ǅ����    �E������������+M;M��  ǅt���    ������������������������+�=�  sz������+U;Usl������f�f����������������������������
u�   ������f�
��������������������f������f����������������q���j j hU  ��x���Q������������++���P������Pj h��  �ؒ��t�����t��� u����E��   �   ǅp���    j �M�Q��t���+�p���R��p�����x���Q�U���E������ x�R����t��p���E���p��������E����t���;�p������t���;�p���~�������+E�E��U����Jj �M�Q�UR�EP�M���U������ x�Q����t�E�    �U��U��	����E�}� ��   �}� t0�}�u������ 	   ������M���U�R����������V�L�E���M������ x�D
��@t�M���u3��%������    �����     ������E�+E�M�3��Q�����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E��t]�����������������̋�U��Qj��������tP�l������E��MQ���������tj�
�����E���]�����������������������������̋�U��} th,Vj jWh�Uj�[�������u�j �������]���������������������������̋�U���tP�������]�����������̋�U��Q��tP�������E��}� t�MQ�U�����u3���   ��]������������������������̋�U��j�h�+h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    �E;�ww9j�������E�    �MQ�������E��E������   �j�����ËE�M�d�    Y_^[��]����������������������������������������������̋�U��Q�E�    �}�wC�EP�������E��}� t�*�=�t u�Y����    ��MQ�H������u����UR�2�����*����    3���}� u�����    �E���]���������������������������������������̋�U����=�t u�����j������h�   �������=�wu,�} t�E�E���E�   �M�Qj ��tR����P�#�=�wu�EP��������E��}� t�E��+�} u�E   �M������M�URj ��tP�����]������������������������������������������������������������̋�U��j�h�+h"�d�    P���SVW�XD1E�3�P�E�d�    �} t�}t	�E�    ��E�   �EԉE܃}� uh@\j jah�[j���������u̃}� u.�n����    j jah�[h|Vh@\�����������b  3҃} �U؃}� uhd[j jbh�[j��������u̃}� u.�
����    j jbh�[h|Vhd[�`����������  j�������E�    �@y�M��	�U�B�E�}� t�M�Q;Uu���}��   �}� th�E�H���U�J�E�H�M��}� uH�U�z t�E�H�U���M�9 t�U��M�Q�P��E�H�@yj�U�R�,������43�uh�Zj jh�[j��������u��E����������    ��   �}� tr�U�B���M�A�U�B�E��M�;@ytM�U�z t�E�H�U���M��E�H�J�U��    �E�@y�H�@y�E��M�@y�h�   h�Zjj褿�����E�}� u�E������S����    �L�U��    �E�@y�H�=@y t�@y�E��M��A   �E�   �U�E�B�M�@y�E������   �j������ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP�,������E��E�    �E���]�����������������̋�U��EP�MQ�UR�EP�MQ�UR�������]���������̋�U��P  ������XD3ŉE��E�    �E�    �} u
�   �  ƅ���� h  ������Pj �0���u8j h<  h�[h�XhXh�!h  ������Q������P�������������U��E�P��������@v]�M�Q�������U��D��E�j hE  h�[h�Xh�`j�xPQ�U�������+й  +�Q�U�R������P�������} t'�EP��������@v�MQ�������U�DÉE��J�����������=����     �}uǅ����xW�
ǅ����L�U���t�M�������
ǅ����L�U���t�}uǅ����dW�
ǅ����L�M���tǅ����t-�
ǅ����L�} t�E�������
ǅ����L�} tǅ����XW�
ǅ����L�} t�M�������
ǅ����L�} tǅ����LW�
ǅ����L�}� t�U��������'�} t�E�������
ǅ����L�������������}� tǅ����H!�
ǅ����L�} tǅ����@W�
ǅ����L������R������P������Q������R������P������Q������R������P������Q������R������P�M�Q�U��lVPh�Vh�  h   ������Q�������D�E�}� }*j h`  h�[h�XhH^j"j�6����R�.����� �&�����������}� }8j he  h�[h�Xh�h��h   ������R�|�����P������h  h�V������P������������������uj�'�����j�����������u�   �3��M�3��w�����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h,h"�d�    P���SVW�XD1E�3�P�E�d�    3��} ���E��}� uhLYj j`h�Xj蒾������u̃}� u-�����    j j`h�Xh�XhLY�j�����3��w  �}�v������    3��_  �=�w��   j�o������E�    �UR��������E܃}� t0�E�    �E;�ww�MQ�UR�E�P�+�������t�M�M��E������   �j�.�����Ã}� uQ�} u�E   �U������U�EP�MQj��tR����E�}� u���P�������������0�   �E������} u�E   �EPj ��tQ����E؋UR�EPj��tQ����E�}� u:�}� @  w�U;U�w��   ��t�E�E�����P�z��������z����0�E�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E������=�t u;h�Y���E��}� thpY�E�P��P��������t��t   ����9�tt4j j�M�Qj ��tR��tP�k������Ѕ�t�}�u	�E�   ��E�    �E��]����������������������������������������������̋�U��j�h8,h"�d�    P���SVW�XD1E�3�P�E�d�    �E�E��} u�MQ��������8  �} u�UR�������3��  �=�w�]  �E�    �}���  j�#������E�    �EP�������E؃}� �  �M;�w��   �UR�EP�M�Q���������t�U�U��j�EP��������E�}� tU�M�Q����U܋E�;Es�M܉M���U�UԋE�P�MQ�U�R�������EP��������E؋MQ�U�R��������}� u{�} u�E   �E������E�MQj ��tR����E�}� tF�E�H����M܋U�;Us�E܉E���M�MЋU�R�EP�M�Q�-������UR�E�P�c������E������   �j�������Ã}� u3�} u�E   �M������M�UR�EPj ��tQ����E���UR�������������    3��K  �}� u	�=�t u;�}� t�+�}� u���P�������������0������    �E��  �EP�r�������u2�}� u���P�O��������O����0��F����    3��   �����   �E�    �}�w(�} u�E   �MQ�URj ��tP����E���MQ�������������    3��e�}� u	�=�t u%�}� t����P�������������0�E��1�UR��������u���P�������������03���K����M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�hX,h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    �} u��   �=�w��   j�ط�����E�    �EP�A������E��}� t�MQ�U�R�&������E������   �j������Ã}� u4�EPj ��tQ�`��E�}� u���P�������������0�3�URj ��tP�`��E�}� u���P�t��������t����0�M�d�    Y_^[��]�������������������������������������������������������������������������������̋�U��j�hx,h"�d�    P���SVW�XD1E�3�P�E�d�    �E������=�wu:j�w������E�    �Ƕ����}�E������E������   �j�k������j j ��tP�̒��u*�����xu�z���� x   �f���� (   ��E������E�M�d�    Y_^[��]�����������������������������������������������������������������̋�U���5���]����̋�U��=�t uh�Bj j?h�Yj�8�������u̃=�t u3���=�wu��w�3�]�������������������̋�U����=�t uh�Bj jgh�Yj�ճ������u̃=�t u3��L  �=�wuv��  ;M҃��U�uh�Zj jph�Yj茳������u̃}� u-�����    j jph�Yh�Zh�Z�d�����3���   �M��w�   ��   �} u
�   �   �=�w��   �}�  w�UR���������t	�E�   ��E�    �E�E��}� u!h(Zj h�   h�Yj�Ӳ������u̃}� u-�U����    j h�   h�Yh�Zh(Z������3��'�U��w��w   �   ������    3���]�����������������������������������������������������������������������������������������������������������������̋�U����} v�}�w	�E�   ��E�    �E�E��}� u!hl[j h�   h�Yj賱������u̃}� u0�5����    j h�   h�YhH[hl[�������   �w3҃=�t �U��}� u!h�Bj h�   h�Yj�G�������u̃}� u0������    j h�   h�YhH[h�B�������   ��M��N3���]������������������������������������������������������������������������������̋�U���3��} ���E��}� u!h�[j h�   h�Yj�y�������u̃}� u0������    j h�   h�Yh�[h�[�N������   �y3҃=�t �U��}� u!h�Bj h�   h�Yj��������u̃}� u0�����    j h�   h�Yh�[h�B��������   ��M��N�3���]������������������������������������������������������������������̋�U��h@  j ��tP����|w�=|w u3��8�M��w�|w��w��t    �xw    ��w   �   ]����������������������������̋�U����xwk�|w�E��|w�M��U�;U�s%�E��M+H�M�}�   s�E���U����U���3���]���������������������������̋�U����E�M+H�M��U����U��   ��M���M#Au�U���u�E�%�  t	�E�   ��E�    �E��]������������������������̋�U���<�E�H�MԋU�E+B�E��M����M�U�i�  �Eԍ�D  �M؋U���U�E����MċUă�t�Y  �E�EĉE��M���ŰE�H��M�Ũ��  �E������E��}�?v�E�?   �M��U��A;B��   �}� sZ�   ��M����ҋE�M�#T�D�E�MԉT�D�U�U��B,�M�M��A�U�U��B��u�   ��M����ҋE#�M��f�M��� �   ����ҋE�M�#���   �E�Mԉ���   �U�U��B,�M�M��A�U�U��B��u�M��� �   ����ҋE#P�M�Q�U��B�M��Q�P�E��H�U��B�A�M�M̉MċU������Uȃ}�?v�E�?   �E���M  �M�+M�M�U������UЃ}�?v�E�?   �E�E�EċM������Mȃ}�?v�E�?   �U�;U���   �E�M�P;Q��   �}� s[�   ��M����ЋM�U�#D�D�M�UԉD�D�E�EЊH���U�UЈJ�E�E��H��u�   ��M����ҋE#�M��f�MЃ� �   ����ҋE�M�#���   �E�Mԉ���   �U�UЊB,�M�MЈA�U�U��B��u�MЃ� �   ����ҋE#P�M�Q�U�B�M�Q�P�E�H�U�B�A�M�M�U��u�E�;E��  �MȋU؍ʉE܋M�U܋B�A�M�U܉Q�E܋M�H�U�B�M�H�U�E�J;H��   �}� sW�U�U��B�M�MȊQ���M�MȈQ��u�   ��M���E�M��   ��M���E�M�T�D�E�MԉT�D�c�U�U��B�M�MȊQ���M�MȈQ��u�Mȃ� �   ���EP�M�Q�Mȃ� �   ���E�M����   �E�Mԉ���   �U�Eĉ�M�MċUĉQ��E؋���U؉
�E؃8 �`  �=�t �B  ��w����tJ�M�h @  h �  �E�P�d��   ���w���tP��t�Q��t�B��wǄ��       ��t�B�HC����t�B�HC��t�Q�BC��u��t�Q�����t�P��t�y���   h �  j ��t�BP�d���t�QRj ��tP�`��xwk�|w��t��+�Q��t��P��tQ蟱�����xw���xw�E;�tv	�M���M�|w��w�E��t�M��w��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���8V�xwk�|w�E�M������MȋU������Ũ}� }����M���E��E�������E�    �M̃� �����UС�w�E�M�;M�s"�U�E�#�M�U�#Q�t��E���E��֋M�;M���   �|w�U�E�;�ws"�M�U�#�E�M�#H�t��U���U��ӋE�;�w��   �M�;M�s�U�z t��E���E���M�;M�uJ�|w�U�E�;�ws�M�y t��U���U��ߋE�;�wu�����E�}� u3���  �M�Q�d������U�J��U�B�8�u3��  �M��w�U�B�E؋M؋�U�}��t!�E�M؋U�#T�D�E�M؋u�#���   �u3�E�    �U�E؋M�#L�D�U�E؋u�#���   �u�M���M��ԋU�i�  �E؍�D  �M��E�    �U�E؋M�#L�D�M�u�E�    �U�E؋M�#���   �M��}� |�U���U��Ẽ��E���M̋U܋D��E��M��+UȉUԋE������E��}�?~�E�?   �M�;M��  �U��E��J;H��   �}� }Z�   ��M����ҋE�M�#T�D�E�M؉T�D�U�ŮB,�M�M̈A�U�U��B��u�   ��M����ҋE�#�M��f�M̃� �   ����ҋE�M�#���   �E�M؉���   �U�ŮB,�M�M̈A�U�U��B��u�M̃� �   ����ҋE�#P�M�Q�U��B�M��Q�P�E��H�U��B�A�}� �  �M��U܍ʉE��M��U��B�A�M��U��Q�E��M��H�U��B�M��H�U��E��J;H��   �}� }W�U�U��B�M�M��Q���M�M��Q��u�   ��M���E��M��   ��M���E�M�T�D�E�M؉T�D�c�U�U��B�M�M��Q���M�M��Q��u�M��� �   ���E�P�M�Q�M��� �   ���E�M����   �E�M؉���   �}� t�U��Eԉ�M�MԋUԉQ��E�EԉE��Mȃ��U��
�Eȃ��M�MȉA��U܋�M܋���M܉��u �U�;�tu�E�;�wu
��t    �M؋U��E���^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�xw;�wuJ��w��k�Q�|wRj ��tP����E��}� u3���   �M��|w��w����w�xwk�|w�E�h�A  j��tQ����U��B�E��x u3��vjh    h   j ����M��A�U��z u�E��HQj ��tR�`�3��9�E��     �M��A    �U��B�����xw���xw�M��Q������E���]���������������������������������������������������������������������������������̋�U���,�E�H�M��U�B�E��E�    �}� |�M���MԋU؃��U���E�i�  �M���D  �U��E�    �	�E���E�}�?} �M�U�ʉE��M��U��Q�E��M��H�ыU����EP�U�jh   h �  �M�Q�����u����/  �U�� p  �U��E�E���M���   �M��U�;U�w]�E��@�����M�ǁ�  �����U����U��E�� �  �M���   �U��J�E�-   �M��A�U����  �U܋E�� �  돋M���  �M�U���E�P�M�Q�U��E��M�H�U����E�P�M�Q�U��E��M�H�U؋E��D�D    �M؋U�Ǆ��      �E��HC�U��BC�U��BC��u�E�H���U�J�   ��M����ЋM#A�U�B�E؋�]������������������������������������������������������������������������������������������������������������������������������������̋�U���0�E������E�M�Q�U܋E�M+H�M�U����U�E�i�  �M܍�D  �U��E���E��M�����UЋE�EЉE��M���U؋E�;E���  �M؃�u�U�U�9U�~3��1  �E������E��}�?v�E�?   �M��U��A;B��   �}� sZ�   ��M����ҋE�M�#T�D�E�M܉T�D�U�U��B,�M�M��A�U�U��B��u�   ��M����ҋE#�M��f�M��� �   ����ҋE�M�#���   �E�M܉���   �U�U��B,�M�M��A�U�U��B��u�M��� �   ����ҋE#P�M�Q�U��B�M��Q�P�E��H�U��B�A�M�M�+M�M؃}� �>  �U�U�U��E������E��}�?v�E�?   �M��U��ʉE�M��U�B�A�M��U�Q�E�M��H�U��B�M��H�U��E��J;H��   �}� sW�U�U��B�M�M��Q���M�M��Q��u�   ��M���E�M��   ��M���E�M�T�D�E�M܉T�D�c�U�U��B�M�M��Q���M�M��Q��u�M��� �   ���EP�M�Q�M��� �   ���E�M����   �E�M܉���   �U��E؉�M�M؋U؉Q��E���M���U���E�E�P��  �M�;M���  �U���E���M���U�U�J��E�E�E��M�+M�MЋU������Uԃ}�?v�E�?   �E؃��1  �M������M��}�?v�E�?   �U��E��J;H��   �}� sZ�   ��M����ҋE�M�#T�D�E�M܉T�D�U�U��B,�M�M��A�U�U��B��u�   ��M����ҋE#�M��f�M��� �   ����ҋE�M�#���   �E�M܉���   �U�U��B,�M�M��A�U�U��B��u�M��� �   ����ҋE#P�M�Q�U��B�M��Q�P�E��H�U��B�A�M�M؉MЋU������Uԃ}�?v�E�?   �EԋM����U�E��M�Q�P�E��M�H�U�E��B�M��Q�E��B�M��U��A;B��   �}� sW�M�M��Q�E�EԊH���E�EԈH��u�   ��M���E�M��   ��M���E�M�T�D�E�M܉T�D�c�U�U��B�M�MԊQ���M�MԈQ��u�Mԃ� �   ���EP�M�Q�Mԃ� �   ���E�M����   �E�M܉���   �U��EЉ�M�MЋUЉQ��   ��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�=�t �  ��w����tA�E�h @  h �  �U�R�d��   ���w���tA��t�B��t�H��wǄ��       ��t�H�QC����t�H�QC��t�B�HC��u��t�B�����t�A��t�z�ub�=xw~Y��t�HQj ��tR�`��xwk�|w��t��+�P��t��R��tP�T������xw���xw��t    ��]����������������������������������������������������������������������������������̋�U���l  �=|w u�����  �|w�E�ǅ����    ���������������������;xw��  �EȋH�M��}� u
������{  �UȋB�E��M���D  �M��UȋB�������E�    �E�    �E�    �	�M���M�}� �  �E�    �E�    �E�    ǅ����    ���������������������@}������Ǆ�����    �Ճ����� �X  �}� u
�������  �M��M��E�    �	�U���U�}��&  �E؃��E܋M܁��  �MЋU܃z��u�EЃ8�t
������u  �M܋�UċEĉ�������������t'�Uă��Uā}�   ~
������=  �E���E��?�M�����������������?~
ǅ����?   �����������������������������}�|�Uă�u	�}��  ~
�������  �E�EċH�;�����t
������  �U�UĉU܋E�;E��-����M�;M�t
������  �U؁�   �U�������E��;M�t
������k  �U��U�ǅ����    ���������������������@��  �E�    �M��M܋U܋B�E��M�;M���   �������E�;��������   �M�;M�r�U��� �  9U�r
�������  �E�% ����E��M����MԋUԁ��  �U��E�;E�t�M�;M�u��Uԋ���EԉE��ދM�;M�u
������  �U������������������?~
ǅ����?   ������;�����t
������U  �U��B;E�t
������@  �M��M܋U����U�������}� t]������ }(�   ���������E�E��   ���������ỦU��,�������� �   ���E��E��������� �   ���U��U��E܋H;M�u�������E�;������t
������   �M��Q;U�t
������   �E����E��&����M�U��E�;D�Du�M�U��E�;���   t������W�M��� �  �M��U���  �U���������������������MȋU�;u�EȋM�;Ht�������Uȃ��U��M���3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h�,h"�d�    P���SVW�XD1E�3�P�E�d�    �L����E��E��Hp#�Vt�U��zl ��   j褎�����E�    �E��Hh�M�U�;�TtI�}� t%�E�P�\���u�}�Ptj�M�Q觚�����UࡨT�Bh��T�M�U�R�X��E������   �j�K�������	�E��Hh�M�}� u
j �2������E�M�d�    Y_^[��]��������������������������������������������������������������������̋�U��j�h�,h"�d�    P���SVW�XD1E�3�P�E�d�    �E�����������E��v����E܋Hh�M��UR��  ���E�E��M;H�  hQ  h�[jh   跅�����E��}� ��  �U܋rh��   �}��E��     �M�Q�UR�y������E؃}� ��  �E܋HhQ�\���u�U܁zh�Ptj�E܋HhQ�������U܋E��Bh�M܋QhR�X��E܋Hp���-  ��V���  j�~������E�    �E��H� u�U��B�u�M��Q�u�E�    �	�E���E�}�}�M�U�E�f�TPf�M�t���E�    �	�E���E�}�  }�M�M�U�A���R���E�    �	�M���M�}�   }�U�U�E䊊  ���S�׋�TR�\���u�=�T�Ptj��TP�ߗ�����M���T�U�R�X��E������   �j��������(�}��u"�}��Ptj�E�P蔗����蔨���    ��E�    �E؋M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h��d�    P��$�XD3�P�E�d�    �E�    �E�P�M�������E�    ��t    �}�u)��t   ����E��E������M�� ����E��}�c�}�u)��t   ����E��E������M������E��N�4�}�u.��t   �M��އ����Q�U��E������M�軧���E���E�E��E������M�衧���EЋM�d�    Y��]����������������������������������������������������������������������������̋�U���,�XD3ŉE�V�EP�������E�} u�MQ�  ��3���  �E�    �	�U����U��}��E  �E�k�0���T;M�+  �E�    �	�U����U��}�  s�EE��@ ���E�    �	�M����M��}�s{�U�k�0�E�����T�M��	�U���U�E����tN�U��B��tC�M���U��	�E����E��M��Q9U�w!�E����T�UU��B��MM��A����v����U�E�B�M�A   �U�BP��  ���M�A�E�    �	�U����U��}�s�E�k�0�M��U�u�f��p�Tf�DJ�ӋMQ�C  ��3��  �����} t!�}��  t�}��  t�UR�����u����k  �E�P�MQ������9  �E�    �	�U����U��}�  s�EE��@ ��M�U�Q�E�@    �}���   �MމM��	�Uԃ��UԋE����tE�U��B��t:�M���U��	�E����E��M��Q9U�w�EE��H���UU��J����E�   �	�E����E��}��   s�MM��Q���EE��P�֋M�QR�\  ���M�A�U�B   �
�E�@    �E�    �	�M����M��}�s3ҋE��Mf�TA��UR�  ��3���=�t t�EP�  ��3�����^�M�3�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M���  �M��}�w-�U�����$���  ��  ��  �	�  �3���]ÍI ���� ������������������������������������̋�U��Q�E�    �	�E����E��}�  }�MM��A ��U�B    �E�@    �M�A    �E�    �	�U����U��}�}3��M��Uf�DJ���E�    �	�E����E��}�  }�MM��U����P�A���E�    �	�M����M��}�   }�UU��E����Q��  �׋�]���������������������������������������������������������̋�U���(  �XD3ŉE�������P�M�QR������-  ǅ����    ���������������������   s��������������������ƅ���� ������������������������������������tD�����������������������������������Q9�����w������Ƅ���� ���j �M�QR�E�HQ������Rh   ������Pjj ������ j �M�QRh   ������Ph   ������Qh   �U�BPj �޸����$j �M�QRh   ������Ph   ������Qh   �U�BPj 觸����$ǅ����    ���������������������   ��   ��������U������t:�M������Q���E������P�M�������������������  �]��������M������t:�E������H�� �U������J�E�������������������  ��E�����ƀ   �2�����   ǅ����    ���������������������   ��   ������Ar?������Zw6�U������B���M������A�������� �E�������  �X������ar?������zw6�M������Q�� �E������P�������� �U�������  ��E�����ƀ   �<����M�3��U�����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�P�M������M��L}���H�y t �M��;}���P�B�E�M������E����E�    �M������E���M��������]������������������������������������̋�U��=$y uj���������$y   3�]����������̋�U��Pw]����̋�U��`w]����̋�U��Q�E���    ��   �M���   �\��   �U���    ��   �E���   �9 ��   �U���    t4�E���   �9 u&j�U���   P�3������M���   R�_������E���    t4�M���   �: u&j�E���   Q�������U���   P������j�M���   R�͉����j�E���   Q蹉�����U���    to�E���   �9 uaj�U���   -�   P膉����j�M���   ��   R�l�����j�E���   ��   Q�R�����j�U���   P�>������M���    \t8�U���   ���    u&�M���   R�)�����j�E���   Q��������E�    �	�U����U��}���   �E����M�|H�Vt:�U����E�|P t*�M����U�D
P�8 uj�M����U�D
PP莈�����M����U�|
L t�E����M�|T uA�U����E�|L u�M����U�|
T t!h�]j h�   hx]j�z������u̋M����U�|
L t:�E����M�|T t*�U����E�LT�9 uj�U����E�LTQ�����������j�UR�Ї������]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�EP�X��M���    t�U���   P�X��M���    t�U���   P�X��M���    t�U���   P�X��M���    t�U���   P�X��E�    �	�M����M��}�m�U����E�|H�Vt$�M����U�|
P t�E����M�TPR�X��E����M�|L t$�U����E�|T t�M����U�D
TP�X�넋M���   �´   R�X���]���������������������������������������������������������������������������������̋�U��Q�} �  �EP�\��M���    t�U���   P�\��M���    t�U���   P�\��M���    t�U���   P�\��M���    t�U���   P�\��E�    �	�M����M��}�m�U����E�|H�Vt$�M����U�|
P t�E����M�TPR�\��E����M�|L t$�U����E�|T t�M����U�D
TP�\�넋M���   �´   R�\��E��]������������������������������������������������������������������������������������̋�U��j�h-h"�d�    P���SVW�XD1E�3�P�E�d�    �����E��E��Hp#�Vt	�U��zl uDj�xw�����E�    ��WP�M���lQ�   ���E��E������   �j�d�������蹨���Pl�U�}� u
j �I������E�M�d�    Y_^[��]�����������������������������������������������������������̋�U��Q�} t�} u3��\�E��M��U�;UtI�E�M��UR�ϋ�����}� t�E�P�������}� t�M��9 u�}��Vt�U�R�|������E��]������������������������������������������̋�U���覧���E��E��Hp����Ƀ��M��U�U��E����E��}�wC�M��$��U��Bp���M��Ap�   �U��Bp����M��Ap�   �   ��V�����u3�t	�E�   ��E�    �E�E�}� u!h`j h�  hx]j�8t������u̃}� u.躒���    j h�  hx]h�_h`�����������E���]Ð��bv�����������������������������������������������������������������������̋�U��j�h(-h"�d�    P��SVW�XD1E�3�P�E�d�    �=�W�VtAj�t�����E�    h�Vh�W��������W�E������   �j舫����ËM�d�    Y_^[��]�����������������������������������������������̋�U��j�hH-h"�d�    P��SVW�XD1E�3�P�E�d�    �} ��   j��s�����E�    �E�x t.�M�QR�\���u�E�x�Ptj�M�QR�������E������   �j說����ËE�8 tcj�ts�����E�   �M�R�������E�8 t#�M��: u�E�8�Vt�M�R�L������E������   �j�?�����ËE� 𭺋M�A�j�UR�C�����M�d�    Y_^[��]�������������������������������������������������������������������������������������̋�U��EP��r����]�������������̋�U��Q�E�    �} |�}�} u3��  hl  h�`jjj�#������E��}� u�u����    3��}  hq  h�`jjh�   �������M���U��: u j�E�P�-~�����-����    3��5  hw  h�`jjh   襍�����M��A�U��z u0j�E��Q��}����j�U�R��}�����ӎ���    3���   h�V�E��Q�E  ���UR�EP�M��R��  ����u3�E��Q�Ǉ�����U��P�G�����j�M�Q�j}�����E�    �x�U��BP�M���BP�q������tDj�M��QR�4}�����E��Q�g������U��P������j�M�Q�
}�����E�    ��U��B�    �M��Q�   �E���]����������������������������������������������������������������������������������������������������������������������̋�U��VW�} t0�} t*�E;Et"�u�6   �}�M�    �UR������_^]�������������������������������̋�U��EP�MQ�e�����]���������̋�U��j�hx-h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    �����E�h�  h�`jjj�8������E�}� u芌���    3��   �|���.����E�M��Ql��E�M��Qh�Pj�o�����E�    �E�Q�%������E������   �j��������j��n�����E�   �U�BP�X��E������   �j�å����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������̋�U���~���]����̋�U��j�h�-h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    �E�    �} |�}	�E�   ��E�    �EԉE؃}� u!h�`j h-  hx]j�kl������u̃}� u0�����    j h-  hx]h�`h�`�@�����3��  �����E���z���U܋Bp���M܉Ap�E�    h8  h�`jjh�   �$������E�}� �8  j�m�����E�   �U܋BlP�M�Q��������E�    �   �j������Ã}� ��   �UR�EP�M�Q�^  ���E��}� ��   �} th�V�UR�`�������t
�u   j�l�����E�   �E�P�M܃�lQ�������U�R��������E܋Hp��u=��V��u2�E܋HlQh�W�r�����j��W��Rhu�]t�����  �E�    �   �j�/��������E�P臂�����M�Q�	������E������   ��U܋Bp���M܉ApËE��M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�졐W�H�0u��W�B�4u��W���   ��W��W���   ��\��W���   �]��W���   ��[��W���   �$]]��������������������������������������̋�U���   �XD3ŉE��} tC�} t�EP�MQ�UR�  ����T�����E���M�TH��T�����T����E��|  ǅd���   ǅh���    �} �O  �M���L�'  �E�H��C�  �U�B��_�  �M��`���hb��`���R�A`������\�����\��� t"��\���+�`�����X���t��\������;u3���  ǅl���   ���l�������l�����l���N��X���Q��`���R��l���k����\Q��y������u"��l���k����\P葔����9�X���u�뚋�\�������\���hb��\���R�^������X�����X��� u��\������;t3��$  ��l���|j h�  hx]h�ahHa��X���R��\���Ph�   ��p���Q��d����P��q������X���Ƅp��� ��p���P��l���Q�UR��  ����t��h�������h�����\����X�����`�����`������t��`�������`�����`�������7�����h��� t�MQ��  ����P����
ǅP���    ��P����U��  �EPj j h�   ��p���Q�UR��~�����E��}� ��   ǅl���    ���l�������l�����l���|��l��� tn��l������U�D
HP��p���Q���������t;��p���R��l���P�MQ�  ����t��h�������h����
ǅd���    ���h�������h����l�����d��� t�MQ��  ���E��0��h��� t�UR�  ����L����
ǅL���    ��L����E���MQ�  ���E��E��M�3��ƈ����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  �XD3ŉE�ǅX���    ǅT���    �Ֆ����D�����D����  ��l���ǅH���   �MQ��@���R��L���Ph�   ��p���Q�UR�\|������u3��  �E���M�THR��p���P蘐������u�M���U�D
H�a  ��p���P�A���������T���h   h�`j��T���Q�#]������X�����X��� u3��  �U���E�LH��8����U�E�L���<���j�Uk��E�L$Q��0���R�ul�����E�H��\���j h  hx]h�bhb��p���R��T�����P��X�����Q�݂����P�lm������X������E���M�TH��L����E�M�T�j��L���R�Ek��M�T$R��k�����}�
  �E��@����H��H�����l����L���T����(�����,���ǅ`���    ���`�������`�����`���;�H�����   �U��`�����l����R;�uJ��`��� t=��`�����l������D���l�����A��`�����l�����(����Ћ�,����L��]�V��`�����l����ЋT���d�����h�����`�����l�����(�������,����T���d�����(�����h�����,����#�����`���;�H�����   j�E�HQ�U�BP��8���Qjh�\jj ������ ����   ǅ$���    ���$�������$�����$���s$��$�����E8������  ��$���f��U8�����h�   ��VP��8���Q�j������u��l����B   ���l����@    ���l����A    ��l����E�H�
�U��l����H���   �}u�U��@����B�MQ�Uk����\�Ѓ���tG�M���U��8����D
Hj��X���Q�m�����U�E��<����L��U��\����B3��   ��8����Vt{�M���U�D
PP�\���uc3�uj j hd  hx]j�_������u�j�E���M�TPR�m����j�E���M�TTR��l�����E���M�DL    ��X��� t��X����   �E���M��X����TP�E���M�DH�M�3�蛂����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�   �E�    �E�    �E�    �E�    �E�U  h}  h�`j�E�P�SW�����E�}� u3��  �M���M��U���U��E��  �M��   �E�   �	�U����U��E����M�THRh8c�E�k����\Qj�U�R�E�P�5U�����}�}kj h�  hx]hch�bhb�M�Q�U�R�(T����P�g�����E������M�THR�E����M�THR詉������t�E�    �  �}� ��   �E�xP tD�M�QPR�\���u33�uj j h�  hx]j�^\������u�j�U�BPP��i�����M�yT tD�U�BTP�\���u33�uj j h�  hx]j�\������u�j�E�HTQ�i�����U�BT    �E�@L    �M�U�QP�E�M��HH�E���   ��   j�U�R�Gi�����E�xP tD�M�QPR�\���u33�uj j h�  hx]j�[������u�j�U�BPP��h�����M�yT tD�U�BTP�\���u33�uj j h�  hx]j�6[������u�j�E�HTQ�h�����U�BT    �E�@L    �M�AP    �U�BH    �E�@h�������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����   �XD3ŉE��Ɍ���   �E�E��(�E��M�� �M�U��,�U��E�   �E��   �E��E��   �E�    �} u3��-  �} t�} u3��  �M���Cuv�E�H��ukj h�  hx]h�dh@dh<d�UR�EP�y����P�d�����} t3ɋUf�
3��Mf�A3ҋEf�P�} t	�M�    �E�  �UR�݅�����E��}��   s0�EP�M�Q���������  �UR�E�P�ۅ��������   ǅ@���    ǅD���    �MQ��H���R�PZ������t3��  ��H���P�M�Q��H���R躄������u3���   �E��H�U��
��H���P�M�Q�U�R��\�����E���t�}��   s�U��@����E���D����
ǅ@���Lj h  hx]h�dh�c��D�����Q��@���R�E�P�M�Q�U����P�b�����} tj�U�R�EP�Na�����} tj�M�Q�UR�6a����j h  hx]h�dh@c�E�P�MQ�UR�w����P�Hb�����E��M�3���z����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��3�]�������̋�U����E�E��E�    �	�M����M��U�;U}A�E����E�j h   hx]hlfh�d�M��Q�R�EP�MQ�M����P�a������E�    ��]��������������������������������������������̋�U���h�   j �EP�������M���u3���  �E���.uX�U�B��tMj h3  hx]hhjhhij�M��Qj�U�   R�eS����P�^`�����Eƀ�    3��e  �E�    �	�M����M�hdi�UR�L�����E��}� u����1  �EE���M��}� uI�}�@sC�U���.t:j hA  hx]hhjhph�E�P�MQj@�UR��R����P��_�����   �}�uI�}�@sC�E���_t:j hD  hx]hhjh�g�M�Q�URj@�E��@P�yR����P�r_�����_�}�uT�}�sN�M���t	�U���,u=j hG  hx]hhjh�f�E�P�MQj�U�   R�R����P�_���������)�E���,u��M���u��U��E�L�M����3���]����������������������������������������������������������������������������������������������������������������������������������������̋�U��j h]  hx]hkh�j�EP�MQ�UR�s����P�$^�����E�H@��t�U��@Rh�jj�EP�MQ�cK�����U���   ��t!�M���   Qh�jj�UR�EP�4K����]����������������������������������������������̋�U���8�EԉE�3Ƀ} ���MЃ}� uhmj jihPkj�R������u̃}� u.�(q���    j jihPkh8khm�~f��������   3��} ���Ẽ}� uh\lj jnhPkj�BR������u̃}� u.��p���    j jnhPkh8kh\l�f��������   �U�U��E��@����M��AB   �U�E�B�M�U��E�Pj �MQ�U�R�������E��} u�E��M�E�H���U�J�E�x |!�M�� 3�%�   �EȋM����E���M�Qj �!f�����EȋE���]����������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�r������]������������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�i������]����������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�ei������]��������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�UR��G������]������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�EP�G������]����������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�h������]����������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�yh������]��������������������̋�U��Q�E�E��M�Q�UR�b������]����������������̋�U��Q�E�E��M�Q�UR�I������]����������������̋�U��Q�E�E��M�Q�UR�EP�}I������]������������̋�U��Q�E�E��M�Q�UR�EP�Y[������]������������̋�U��E��=   vh@lj j8h�kj�TN������u̋UR�EPj ��G����]����������������������������̋�U����EP�M��X���M����   vh@lj jDh�kj��M������u̃}�|5�}�   ,�M��8M��� ���   �U�Q#E�E�M��m���E��1�'�M��M������   �B�#E�E�M���l���E���M���l����]��������������������������������������������������̋�U���(�EP�M��1W���}�|6�}�   -�M��L������   �E�B#M�M��M��[l���E��   �M��WL��P�U�����   R�QN������t!�E��%�   �E�M�M��E� �E�   ��U�U��E� �E�   j�M��L��� �HQ�M���K����BP�M�Q�U�R�E�Pj�M���K��P�S����� ��u�E�    �M��k���E���M�#M�M؍M��k���E؋�]������������������������������������������������������������������������������̋�U��=u u�E��W�A#E��j �UR�EP�*b����]��������������������������̋�U��E�U��DV�u�     j�E�P3�NVf�
�����u3�^��]ËM�U�E�QRP�����t�U��MZ  f9
u֋B<��~�8PE  u��HSW�x�D+�3�3ۅ�v���;�r	��+�;p�rC��(;�r�;�t[C�=Du u �=@u uH�  �@u��t:�Du��@uh�lP��3�;�t�U�R�UVV�M�QVVVR�Ѓ� ��u	_[3�^��]ËM����u���=��1��  �M���@�U�Rh�lV�Ѕ��u  �M��R VVV�E�PWS�҅��P  �M�u���@h�U�R�Є��-  �M�;��"  ��B�Ѕ���   �M���Rj �E�P�E�P�EP�E�Pj �҄���   �E;�u�E�;�w	�M��;�r�M���B�Ѕ�u��   �E�����   =�����   ��    Qj ���P���������   �M���RV�E�Pj j j �E�P�҄�tU+}�;>rN�M��   ;�v�I ;<�r@;�r��D���Mj %��� ��M��Rpj j �EP�EP�E�P�҄�t�E�   Vj ���P�`��M����ҋM��P@�ҋM��P8�ҋM���P(�ҋE�_[^��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  �XD3ŉE��=Hu t3��M�3��sk����]á�WV�5�P�Hu   �օ��x  h,m�֋���u^�M�3��6k����]�S��hmV�Ӊ�������u[^�M�3��k����]�WhmV�Ӌ����  h�lV�Ӌ؅��
  ������Qjj h�lh  �����������   ������������RP������Pj h�lQ�ׅ���   ����������+Ѓ���   ��=  ��   ������P������������Q������Rj h�lP�׋�����Q����V�����ua�������\8�����t	�������I�������5�W3���������@��~�����P��_[^�M�3���i����]�V���_3�[�M�3�^��i����]��������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��Q�E�   �} u�E�    �E���]������������U��SVWUj j h�C�u�({��]_^[��]ËL$�A   �   t2�D$�H�3��h��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h�Cd�5    �XD3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y�Cu�Q�R9Qu�   �SQ��W�SQ��W�L$�K�C�kUQPXY]Y[� �������������������������������������������������������������������������������̋�U����E%�����E�M#M��������   �} tj j �El�����U�3�t	�E�   ��E�    �M��M��}� uh�mj j1h`mj�JC������u̃}� u-��a���    j j1h`mh<mh�m�"W�����   �/�} t�EP�MQ�k�����U���EP�MQ�k����3���]����������������������������������������������������������������̋�U����EP�M��L���M���A����t2�M���A������   ~�M���A��Ph  �UR��X�����E��h  �EP�M��A��P��;�����E�M�M�M��a���E��]��������������������������������������������̋�U��=u uh  �EP�i>������j �MQ�_O����]�������������̋�U����EP�M��K���M��A����t/�M���@������   ~�M���@��Pj�UR��W�����E��j�EP�M���@��P��:�����E�M�M�M��`���E��]����������������������������������̋�U��=u uj�EP�=������j �MQ�dl����]����������������̋�U����EP�M���J���M��#@����t/�M��@������   ~�M��@��Pj�UR�W�����E��j�EP�M���?��P�:�����E�M�M�M��_���E��]����������������������������������̋�U��=u uj�EP�<������j �MQ��Q����]����������������̋�U����EP�M���I���M��C?����t/�M��7?������   ~�M��$?��Pj�UR�$V�����E��j�EP�M��?��P�49�����E�M�M�M���^���E��]����������������������������������̋�U��=u uj�EP��;������j �MQ�JL����]����������������̋�U����EP�M��I���M��c>����t2�M��W>������   ~�M��D>��Ph�   �UR�AU�����E��h�   �EP�M��>��P�N8�����E�M�M�M���]���E��]��������������������������������������������̋�U��=u uh�   �EP��:������j �MQ��E����]�������������̋�U����EP�M��H���M��s=����t/�M��g=������   ~�M��T=��Pj�UR�TT�����E��j�EP�M��2=��P�d7�����E�M�M�M��]���E��]����������������������������������̋�U��=u uj�EP��9������j �MQ�bb����]����������������̋�U����EP�M��1G���M��<����t/�M��<������   ~�M��t<��Pj�UR�tS�����E��j�EP�M��R<��P�6�����E�M�M�M��,\���E��]����������������������������������̋�U��=u uj�EP�9������j �MQ��P����]����������������̋�U����EP�M��QF���M��;����t2�M��;������   ~�M��;��Ph  �UR�R�����E��h  �EP�M��l;��P�5�����E�M�M�M��F[���E��]��������������������������������������������̋�U��=u uh  �EP�)8������j �MQ��Q����]�������������̋�U����EP�M��aE���M���:����t2�M��:������   ~�M��:��PhW  �UR�Q�����E��hW  �EP�M��|:��P�4�����E�M�M�M��VZ���E��]��������������������������������������������̋�U��=u uhW  �EP�97������j �MQ��N����]�������������̋�U����EP�M��qD���M���9����t2�M���9������   ~�M��9��Ph  �UR�P�����E��h  �EP�M��9��P�3�����E�M�M�M��fY���E��]��������������������������������������������̋�U��=u uh  �EP�I6������j �MQ��d����]�������������̋�U����EP�M��C���M���8����t/�M���8������   ~�M���8��Pj �UR��O�����E��j �EP�M��8��P��2�����E�M�M�M��|X���E��]����������������������������������̋�U��=u uj �EP�l5������j �MQ�FN����]����������������̋�U��}�   ���]��������������̋�U��E��]���̋�U��Q�EP�MQ�
F������u�}_t	�E�    ��E�   �E���]�������������������������̋�U��Q�EP��6������u�}_t	�E�    ��E�   �E���]�������������̋�U��Q�EP�MQ�NN������u�}_t	�E�    ��E�   �E���]�������������������������̋�U��Q�EP�7������u�M��_t	�E�    ��E�   �E���]�������������������������̋�U��E�� ]���̋�U���4�EP�M��1A���}   ��   �M��6����t/�M��z6������   ~�M��g6��Pj�UR�gM�����E��j�EP�M��E6��P�w0�����Ẽ}� t,�M��+6������   �E��M��M��V���E��*  ��U�U܍M���U���E��  �M���5��� ���   ~D�M���5��P�M�����   Q��7������t"�U�����   �U��E�E��E� �E�   ��T��� *   �M�M��E� �E�   j�M��t5����BPj�M�Q�U�R�E�Ph   �M��S5����QR�M��E5��P��m����$�E�}� u�E�E؍M��U���E��A�}�u�M��MԍM���T���E��'��U��E���ЉUЍM���T���E���M���T����]����������������������������������������������������������������������������������������������������������������������������̋�U��Q�=u u$�}A|�}Z�E�� �E���M�M��E���j �UR�h`������]���������������������������̋�U���@�XD3ŉE��E�    �E�    �EP�M��i>���M���3��Pj j j j �MQ�U�R�E�P�G���� �E��MQ�U�R�}T�����E��E���u8�}�u�E�   �M��oS���E��j��}�u�E�   �M��SS���E��N�:�M���t�E�   �M��5S���E��0��U���t�E�   �M��S���E���E�    �M��S���E��M�3��W����]�������������������������������������������������������������������������������̋�U��j �EP�MQ��_����]�������̋�U���@�XD3ŉE��E�    �E�    �EP�M���<���M��[2��Pj j j j�MQ�U�R�E�P�2F���� �E��MQ�U�R�k�����E��E���u8�}�u�E�   �M���Q���E��j��}�u�E�   �M���Q���E��N�:�M���t�E�   �M���Q���E��0��U���t�E�   �M��Q���E���E�    �M��Q���E��M�3��U����]�������������������������������������������������������������������������������̋�U��j �EP�MQ�d����]�������̋�U���@�XD3ŉE��E�    �E�    �EP�M��;���M���0��Pj j j j �MQ�U�R�E�P��D���� �E��MQ�U�R��Q�����E��E���u8�}�u�E�   �M��P���E��j��}�u�E�   �M��sP���E��N�:�M���t�E�   �M��UP���E��0��U���t�E�   �M��7P���E���E�    �M��#P���E��M�3��0T����]�������������������������������������������������������������������������������̋�U��j �EP�MQ�d����]�������̋�U����E�E��M�Q�U�3��} ���E�}� uht�j j7h�nj��/������u̃}� u0�N���    j j7h�nh�nht���C�����   �$  3�;U��؉E�uh��j j8h�nj�/������u̃}� u0�N���    j j8h�nh�nh���sC�����   ��  �U� 3��} ����#E��;E��ىM�uhPnj j=h�nj�#/������u̃}� u0�M��� "   j j=h�nh�nhPn��B�����"   �J  3��} ���E�}� uh0nj j>h�nj�.������u̃}� u0�?M���    j j>h�nh�nh0n�B�����   ��   �U��0�E����E��} ~A�M����t�E���M�U����U���E�0   �E��M��U����U��E���E빋M�� �} |>�U����5|3�M����M��U����9u�M��0�U����U���E�����U��
�E���1u�U�B���M�A�&�U��R�Z������P�E��P�MQ�6����3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���,�XD3ŉE��EP�M�Q�_�����U�Rj j���ċMԉ�U؉Pf�M�f�H�vd�����U�B�E�M��U��E�Pj j.h�oh�ohho�M�Q�UR�EP�L����P�7�����M�U�Q�E�M�3���O����]���������������������������������������������������̋�U����E�   �3�f�E��M�Q���  ��f�U��E�H�� �  f�M�U�B%�� �E�M��U��E��E�}� t�}��  t�P��  f�M��a�}� u)�}� u#�U�B    �E�     �Mf�U�f�Q�   �E�<  f�E��E�    ��M����  f�M��U����?  f�U��E���E��M�����U�B�E����M��U�B%   �u;�M�Q��E���   ������ыE�P�M���E�f�M�f��f�M���U��E�ЋMf�Q��]���������������������������������������������������������������������������������������������̋�U����Lu�E��M�����Ƀ��M�uh0qj j*h�pj�$*������u̃}� u+�H���    j j*h�phxph0q��=�����E���E�Lu�E���]��������������������������������̋�U��Lu]�����SW3��D$�}G�T$���ڃ� �D$�T$�D$�}�T$���ڃ� �D$�T$�u�L$�D$3���D$���3�OyN�S�؋L$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$Oy���؃� _[� ����������������������������������������������WVS3��D$�}G�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u�L$�D$3���؋D$����A�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�Ou���؃� [^_� �����������������������������������������������������̀�@s�� s����Ë�3������3�3������������������̀�@s�� s����Ë�3Ҁ����3�3�������������������U��W�}3�������ك��E���8t3�����_��������������������̋�U��j�>����]���������������̋�U��j�h�-h"�d�    P�ĘSVW�XD1E�3�P�E�d�    �} u3��   j��"������u3��oj�(�����E�    �EP�MQ�Pu�Y���URj �EP�MQ�UR�M��LD���M��kE���E�Pu�Q���E������   �j��^����ËE�M�d�    Y_^[��]��������������������������������������������������������������̋�U��Q�M��E��M��U��E�B�M��A    �U��B    �E��@    ��]� �����������������̋�U��Q�M��E��x t7�M��U��B�A�M��y t"�U��B�M���Q�E��HQ�U��B�Ѓ��ɋ�]�������������������̋�U��j�h.h"�d�    P�ĘSVW�XD1E�3�P�E�d�    �} u3��   j�!������u3��pj�X&�����E�    �EP�MQ�Pu��W���U R�EP�MQ�UR�EP�M��B���M��C���E�Pu��O���E������   �j�]����ËE�M�d�    Y_^[��]�������������������������������������������������������������̋�U��Q�M��M��JB���M���,�?B���E�tu�tu�pu�} t�U�|u�E�xu��xu    �|u    �M���,�hu�U��du�E��u�M��u��u �E���]� ��������������������������������������������̋�U���H�M��M��jP���M��bP���=tu ��   �tu���?uG�tu�B��@u8�pu���pu�U�R�)����Ph�y�E�P��1����P�M��
���v�tu���?uS�tu�H��$uEj �U�R�7����P�M������M��L����u�tu�pu�M�Q�>)����P�M������U�R�')����P�M�����M��wL����u	3��  �?�M��aL����t�{7����u�pu���t�tuR�M���S����E�P�M��=���=xu u2�M��?�����|ujhPu�|uQ��"�����E��U��xu�=xu ��   �|uP�xuQ�M��3���xu�U�E�E�M����tY�E���� u0�U���U�E��  �M���M�U���� u�M���M�����U�E��
�U���U�E���E�띋M�U���xu��]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�M�jPh�u�M��p2����u��]���������������̋�U���h��-����tH��u%������uj �M�Q�������u��    ��u�E�P�M�,���E�  �  �pu���?�t  �pu���pu�pu���?uK�pu�H��?u=�U�R�&�����pu���t�pu���pu��E�P�M�+���E�9  �M�Q�M�����M��/ ���E�M���%���E��M��(����u�U�R�M�D+���E��  �pu�����   �pu���@��   �M�Q�zD�����M���(������   ��u��tn��u �E�P�M�Q�M��=G��P�M�����pu���@t>�M�Q�%D����P�M������U�R�E�Ph�y�M�Q�M��Q������F��P�M������)�U�R�E�Ph�y�M�Q�M��hQ������F��P�M�����}� t�M���)���}� t�M��t#���M���'����u�M���)����t�U�R�M�*���E��   �   �pu���t�pu���@ut�pu���t�pu���pu�,3����t:�}� u4�M��L$����u(�M���J��P�M�Q�<�����U�R�M�)���E�U��E�P�MQ�d<�����E�>�j�M��V���E�-�+�pu���tj�M�V���E��j�M�V���E��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��pu���?uJ�pu�B��$uj�MQ�51�����E�;�$�pu���puj j �EP��=�����E��j j�MQ�	R�����E]�������������������������������̋�U���h�XD3ŉE�pu���0�M�x5�}�	/�pu���pu�E�P�MQ�hu�g���E�;  �6  �M��H���pu���?ubj �M�Q�Y0����P�M�����pu��pu���pu��@t)�pu���pu�pu�����ك�Q�M��TB���  jh�y�puR��  ����u�E��y�pu���pu�9jh�y�puQ��  ����u�E��y�pu���pu��E�    �}� ��   �E�P�D?������"����twj�M�Q�M��,���U�R�_8����P��u���EЃ}� t�E�P�M��=L���:h�y�M��.L��h�y�M�Q�U�R�E�P�M�Q�A)�������M��P�M��~���:h�y�M���K��h�y�U�R�E�P�M�Q�U�R�)��������L��P�M��B���N�E��t.�pu���@u �M���F��P�M������pu���pu�j@hpu�M��)��P�M������M��t�hu�Q����u�U�R�hu����E�P�M�U%���E�M�3��&=����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  �M��E���M��E���E�    �E�    �pu�������pu���pu���������������_�o  �������lx�$�Px�pu���puj�M�UQ���E�  �M��3E���M����   �U�R�:����Pj<�E�P�I����P�M��0���M��/���ȃ�>u
j �M��g:��j>�M��]:���} t�U��pu���u�U�R�M�}#���E�  �pu���pu�pu�M�j j �U�R�UM����P�M�����Eܣpu�M��� ����u*�pu�Q���1u�E�Pj~�M�Q��H����P�M��M���M�� ����u�U�R�M��[���E�P�M��"���E�v  �%  �pu�Q���hwP�M��H���  �E�   �pu�Q���LwP�M��H����  �pu�������pu���pu���������������_��  ������� y�$��x�pu���puj�M�O���E��  �pu�B����wQ�M���G���F  �pu�B����wQ�M�Q���E�  �  �pu�B����wQ�M��*���M������U�R�M�!���E�F  ��  jhhv�E�P������M��3H���M�Q�M�!���E�  �pu�B����wQ�M�����E��  �pu�B����wQ�M��*G��j j �U�R��6����P�M��h���M�������u�M��bA����tj�M�QN���E�  �E�P�MQ�M��J=���E�{  �  �  �pu�B����wQ�M��F���pu���uj�MQ�M��6���E�4  �pu���0�E�x�}�rj�M��M���E�  �M���xR�M��LF���pu�������pu���pu�����������������0�����������>  ������$�`yj �E�P�������M�Q�UR�E�P��t���Qj ��|���R�M��2;�����4<�����-<���E�^  �  �E�P�M�Q�M��<��j,��d���R��l���P�J8��������:��P�M�����j,��T���Q��\���R�"8��������:��P�M�����j,��D���P��L���Q��7�������:��P�M����j)��4���Rj ��<���P��J�������n:��P�M��x��j'�MQ�M��W:���E�  �;�U�R�EP�M��F;���E�w  �!�pu���puj�M�L���E�T  ��  �pu�B����wQ�M��D����  �pu��� ����pu���pu�� ��������������� t������0t!�N�pu���puj�M�K���E��  j h�y�M�Q������M���D���U�R�M����E�  j�M�PK���E�  �0  �pu��������pu���pu��������������������A������������	��   ��������|y�$�ty�pu�Q���@xP�M�����E�  �pu�Q���@xP�M������pu���?u5��,���P�����P�M�����pu���@u�pu���pu���$���Q�V?����P�M��n��h�y�M��k%���U�R�M�����E��j�M�)J���E�n�j�M�J���E�]�j�M�J���E�L�}� t
�M��J���-�M��V����u!�E�Ph,w�����Q�����P�M��	���U�R�M�i���E��]ÍI �p�p�q�q�qr�w fr�r�r�rv7ssYs�s�s�u�v�w 	

�t�t�u�u�uw7w        �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M�����pu��pu���pu��@u�pu��pu���pu��_tj�M��E���E�   �pu���puj �U�R�#D����j �E�P�D�����pu���t�pu���@t�pu���pu�աpu���u�pu���puj�M�HE���E��pu���pu�M�Q�M�����E��]��������������������������������������������������������������������̋�U����   �M��8���E� �M��5������  �pu�����  �pu���@��  ��u��t��u��u�E�P�M�$���E�(  �M�������uE�M�Qh�y�U�R�����P�M��7���E���t�M�Qj[�U�R�<����P�M�����E� �pu���?�  �pu���pu�pu���@�����@�����$��@�����@���%��  ��@�����Ԁ�$����pu�B��_ua�pu�Q��?uR�pu���pu�M�Q�U�Rj j �E�P��+�������2��P�M��_���pu���@u�pu���pu�@�M�Q�U�Rj'�E�P�M�Q�����Pj`�U�R�;�������%1�����'2��P�M������   �pu���pu�M�Q�U�Rj j�E�P�?��������1��P�M�������   j@hpu�M��z���M�Qh�y�U�R�x����P�M�����hu�#����u�E�P�hu�����w�pu���pu�U�R��|���Pj]�M�Qj j�U�R�?�������R0�����T1��P�M��/���E��*�E�P��l���Q��t���R�)�������$1��P�M������.�E�P��\���Qj j��d���R�>��������0��P�M����������pu���<�����<��� t��<���@tW�W�M������tj�M��/���;�U�R��D���Ph�y��L���Qj��T����xA�����;�����{0��P�M��V����
j�M��B/���U�R�M�����E��]Ð�~1B~~� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����pu���uj�M��?���E�T�R�pu���?u3�pu���puj �U�R�<>����Pj-�EP�88�����E��j �MQ�>�����E��]�������������������������������������̋�U���   V�E�    �pu���Qu�E�z�pu���pu�pu���uj�M�#?���E�S  �N  �pu���0��   �pu���9��   �}� tG�pu� ��/��E��U��pu���pu�U�R�E�P�M��
��P�M�Q�U�R�x�����E��4�pu� ��/��E��U��pu���pu�U�R�E�P�M������E��M��M�U�R�M����E�  �  �E�    �E�    �pu���@��   �pu���uj�M�>���E�L  �W�pu���A|7�pu���P*�E��U�������ȋ�pu���A���M��u��j�M��=���E��   �pu���pu�e����pu��pu���pu��@tj�M�=���E�   �M��tX�}� t&�U�R�E�P�M����P�M�Q�U�R������E���E�P�M�Q�M��i���E��U��UЋE�P�M�����E�V�T�}� t&�M�Q�U�R�M��U��P�E�P�M�Q�������E���U�R�E�P�M��/���E��M��M��U�R�M�{���E^��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����pu���u3���   ��   �pu���0|8�pu���9*�pu���/�M��pu���pu�E��   �   �E�    �pu���@tY�pu���u3��k�7�pu���A|$�pu���P�U����pu��T
��U������2�pu���pu뚋pu��pu���pu��@t�����E���]����������������������������������������������������������������������̋�U����   �pu���?u�pu�B��$tj�M�:���E�  �pu���pu�du�U��hu�E̋lu�M���\����n���M��f���M��^����\����du�E��hu�MЉlu�M��.���M��.���E� �pu���?u/�pu���pu�U�Rj��T���P�_"����P�M�������jj��L���Q�6����P�M������M��,
����t��u�U���up��D���P��"����Pj<��<���Q�2����P�M�� ���M��u���Ѓ�>u
j �M���"��j>�M���"���E��t�pu���t�pu���pu�M��du�Ủhu�E��lu�M�Q�M�����E��]�����������������������������������������������������������������������������������������������������������������̋�U���|�XD3ŉE��E�   �M��l,����u�M��Q)�����  �pu����  �pu���@��  �}� t	�E�    �
j,�M��!���pu���0�U�x4�}�	.�pu���pu�M�Q�U�R�lu�w���P�M������  �pu�E�M���+���pu���Xu�pu���puhTz�M��M0���%  �pu���$u7�pu�H��$t)�pu���pu�E�P�k����P�M��_�����   �pu���?��   �E�P�"�����U����tkj�M�Q�M������U�R������P��u���Eă}� t�E�P�M��/���.h�y�M�Q�U�Rh<z�E�P��������0��P�M�������.h�y�M�Q�U�Rh<z�E�P��������Z0��P�M�������M��*��P�M�Q��$����P�M��z����pu+U��~�lu�������u�E�P�lu�����M�Q�M��h����������u �U�R�M�����E�M�3�� ����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  �XD3ŉE�pu��M��pu���pu�E�������������R��  �����������$����EP�} �����E�  �pu���@u$�pu���puh\z�M������E�S  �3��D���Q�R����P�URhw��L������������#���E�  �EP�"�����E�
  �M�Q�������U�R�������M��m������   �M��]����t{jd�E�P�M������uj�M�I4���E�  �M��M��U���-u�E��E��E�.��E�.�M�Q�URje��4���P�M�Q��<����������"�����#���E�]  �j�M��3���E�I  ��x���R�,����������tSj��h���P��x����e����h���Q�>����P��u����d�����d��� t��d���R�M�����E��  �E���Du5h�y�MQ��x���Rh<z��,���P�	��������,���E�  �3h�y�MQ��x���Rhz��$���P���������,���E�m  �h  j j ��\���Q�/���������R�8������\���P�M�v���E�/  j{��T�����
���M�������������H|3������J~�(�����R� ����P��T�������j,��T��������E���������������F������������wx�������$��������P�����P��T����=���j,��T�����������Q�i����P��T�������j,��T����Y��������R�A����P��T��������j}�EP��T��������E�-�+�pu���puj�M�1���E�j�M�1���E�M�3������]Ë�E�ٌ�f�'�R�A��c� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  �M��#���A���E��M�!����E��}���  uj�M�/���E�  �B�}���  u�EPj�MQ�r,�����E�  ��}���  u�UR�M����E�j  �E�% �  �0  �M��� �  t�U���   3���   ���������M��� `  ��Ƀ����������� t�U���   �� �����E�%   �� ����� ��� t>�M��� �  t�U���   3���   ���������
ǅ����    ������ ��
  �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ t|�M��� �  t�U���   3���   ���������
ǅ����    ������ ��	  �M��� �  t�U���   3���   ���������
ǅ����    ������ ��	  �M��� @  tM������t/�A����t&�U�R�E�����Pj �E�P��%����P�M��Z�����M�Q������P�M������U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� t�E�%   ��������M���   ������������ �-  �U��� �  t�E�%   3�=   ���������
ǅ����    ������ ��   �U�R������P��|���Pj{�M�Q�M��������P�M������U�R�B������e����u1h�{��l���P�M�Qj,��t���R��$��������%��P�M��E���h�{�M��B���E�P������������tR������tI� ����u@�M�Q��T���Rj ��\���P�M�Qj ��d���R�U$����������������P�M������  �M�����M�����M�����M�����M��w���E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t�M���   ��������U���   ������������ �"  �E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t[�M���   ��   uJ��L���R�R����P�M�������D���P�:����P�M�������<���Q�"����P�M��p����k�U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� t'�E�%   =   u��4���Q�����P�M�������,���R�����P�M�������E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� ��   �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t8�U��� �  t�E�%   3�=   ���������
ǅ����   ������ u;�v�����t��$���R�&����P�M�����������P�&����P�M��k��������tO�����t,�M�Q�����R�����P�����������P�M�����������Q�����P�M�����������R�w����P�M������M�������uA�M��������u)�n����u �EPj ������Q�� ����P�M��a�����UR�M��-����E�    �M�����}� tNj ������P�l����Ph ������Q�������P�M�����������t�U�R�M�����E��  �bj hPuj�x����������������� t����������������
ǅ����    �������E��M�Q������R������P�M��h����E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t�M���   ��������U���   ������������ ��  �E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� ��   �M���   ��   uzj,������R�E�P������Qj,������R�E�P������Qj,������R�E�Ph�{������Q�.��������a�����c�����S�����U�����E��P�M��O����   �U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� tB�E�%   =   u3j,������Q�U�Rhp{������P�����������P�M�������h`{�M��� ��h�{������Q�M��4��P�M�����j)��x���R������P�3����Pj(������Q���������V��P�M��`����U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� ��   �E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t:�M��� �  t�U���   3���   ���������
ǅ����   ������ u�M�Q�M������g�����t��p���R�����P�M��m������h���P�����P�M����������t�}� t�M�Q�M������U�R�M������  �EP�M������M��� �  u.�U��� |  �� h  u�E�P�MQ�������E��	  �1  �U��� �  u,�E�% |  = p  u�M�Q�UR�0������E�	  ��  �E�% �  u]�M��� |  �� `  uLh�{�UR��X���P�@�����P��P���Qj{��`���R�M��L�����N���������E�N	  �  �E�% �  u.�M��� |  �� |  u�U�R�EP�������E�	  �[  �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ tL�M��� �  t�U���   3���   ���������
ǅ����    ������ th8{�M��a����  �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ tL�M��� �  t�U���   3���   ���������
ǅ����    ������ th�z�M�������   �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ tI�M��� �  t�U���   3���   ���������
ǅ����    ������ th�z�M�������0�M��� �  u%�U��� |  �� x  u�E�P�M�N����E�  �M��� �  t�U���   3���   ����|�����M��� `  ��Ƀ���|�����|��� t�U���   ��x�����E�%   ��x�����x��� ��   �M��� �  t�U���   3���   ����t����
ǅt���    ��t��� u:�M��� �  t�U���   3���   ����p����
ǅp���    ��p��� t#�M�Qh ��H���R�f�����P�M�������E�P��@���Q�`�����P�M��f����U��� �  t�E�%   3�=   ����l�����U��� `  ��҃���l�����l��� �x  ������R  �E�% �  t�M���   3ҁ�   ��h�����E�% `  �������h�����h��� t[�M��� �  t�U���   3���   ����d����
ǅd���   ��d��� t!�M�Qh�z��8���R�T�����P�M��r����E�% �  t�M���   ��   �s  �U��� �  t�E�%   3�=   ����`�����U��� `  ��҃���`�����`��� t�E�%   ��\�����M���   ��\�����\��� �$  �U��� �  t�E�%   3�=   ����X�����U��� `  ��҃���X�����X��� t�E�%   =   ��   �M��� �  t�U���   3���   ����T�����M��� `  ��Ƀ���T�����T��� t�U���   ��   tU�E�% �  t�M���   3ҁ�   ��P�����E�% `  �������P�����P��� t2�M���   ��   u!�U�Rh�z��0���P������P�M������������  �M��� �  t�U���   3���   ����L�����M��� `  ��Ƀ���L�����L��� tl�U��� �  t�E�%�   3Ƀ�@����H�����U���   3���   ����H�����H��� t&�M�Qh�z��(���R�������P�M������Z  �E�% �  t�M���   3ҁ�   ��D�����E�% `  �������D�����D��� tp�M��� �  t�U����   3����   ����@�����M���   3ҁ�   ��@�����@��� t&�E�Ph�z�� ���Q�3�����P�M��Q����   �U��� �  t�E�%   3�=   ����<�����U��� `  ��҃���<�����<��� tb�E�% �  t�M����   ��Ƀ���8�����U���   ��҃���8�����8��� t!�E�Ph�z�����Q������P�M������U��� �  t�E�%   3�=   ����4�����U��� `  ��҃���4�����4��� t�E�%   ��0�����M���   ��0�����0��� t*�F�����u!�U�Rhtz�����P�������P�M������M���   t!�U�Rhdz�����P�������P�M�������M�Q�M�����E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���x�E�    �pu���_u�U��� @  �U��pu���pu�pu���A�  �pu���Z�  �pu���A�E��pu���pu�U��� �  �U��E���t�M���    �M���U��������U��}���  �E�% �  t�M���������   �M��U��U���E�%�����E��M��M�U����U�t�}�t@�}�tq�   �E�% �  t�M���?�����@�M���U���������   �U��E��E��r�M��� �  t�U���?����ʀ   �U���E�%����   �E܋M܉M��;�U��� �  t�E�%?����E���M��������M؋U؉U���E���  �E��k  �E����Eԃ}���   �M��$����U���������   �U��   �E�%����   �E��s�M��� �  t�U���������   �U��;�E�% �  t�M���������   �M��U��U���E�%�����E��M��M̋ỦUЋEЉE����E���  �E��  �  �pu���$��  �E� �pu���pu�pu��Uȃ}�R�]  �E������$�Զ�U����d���� �  �U��D  �E�%�g�� �  �E��/  �M����d���� �  �M��  �U����d���� �  �U��  �E�%���� |  �E���  �pu�Q��Pu�pu���pu�pu���pu�pu��Eă}�Q��   �M���d��$�P��pu���pu�h����  �pu���pu�pu���0|C�pu���95�pu��pu�D
ѣpu�����E��M���   �M��E��-  ��E���  �7�pu���pu������	  �E���  �E���  �E���  �E���  ��  �E���  �pu���pu��  �E��pu���pu�pu���0|�pu���5~$�pu���t	�E���  ��E���  �E��z  �pu���0�E��M��� �  �M��U��� �  t�E�%����   �E��M��M���U��������U��E��E��M���t�U���������   �U���E�%����   �E��M���t�U���    �U���E�%�����E��M����M�t�}�t@�}�tr�   �U��� �  t�E�%?�����@�E���M���������   �M��U��U��s�E�% �  t�M���?����ɀ   �M���U���������   �U��E��E��;�M��� �  t�U���?����U���E�%�����E��M��M���E���  �E��  ��E���  �E��  �pu���pu��  �pu���0��  �pu���8��  �pu��U�pu���pu�M�������M��U�U��E���0�E��}��?  �M��$����U��� �  t�E�%����   �E��=�M��� �  t�U���������   �U��E��E���M��������M��U��U��E��E��M��M��U��� �  t�E�%?�����@�E���M���������   �M��U��U��  �E�% �  t�M���������   �M��;�U��� �  t�E�%����   �E��M��M���U��������U��E��E��M��M��U��U��E�% �  t�M���?����ɀ   �M���U���������   �U��E��E��  �M��� �  t�U���������   �U��;�E�% �  t�M���������   �M��U��U���E�%�����E��M��M��U��U��E��E��M��� �  t�U���?����U���E�%�����E��M��M��   �U��������� @  �U��l�E�%���� `  �E��Z�M���������    �M��F�U��������� h  �U��2�E�%���� p  �E�� �M��������� x  �M���E���  �E��H�C�pu���9u�pu���pu�E���  ��pu���t	�E���  ��E���  �E���]ÍI �����z��c�˱��7�N�e���z������ 																																																																					����&����� ��(���Z�����#�7�I������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���j �������P�M������pu���tl�pu��E�pu���pu�U�U�}�0t�}�2t�}�5t(�5hTz�M��K����&�E�P������P�M��*����j�M����E�(�
j�M������h�{�M��
����M�Q�M�����E��]���������������������������������������������������̋�U���@�M��}���j j�E�P�5����P�M��k����M��P�����uN�pu���tA�pu���@t4�U�R�E�Ph�y�M�Q�U�R�O���������������6���P�M������pu���@u�pu���pu�b�pu���tj�M�������J�M��J�����tj�M������2�U�R�E�Ph�y�M�Qj�M�������X���������P�M������U�R�M�@����E��]��������������������������������������������������������������������������̋�U����pu����  �pu���A�E��pu���pu�}���   �M��������������   �U�����U��}���   �E�����$��j�0�����P�M��Q����gj������P�M��<����Rj������P�M��'����=j�������P�M������(j�������P�M�������j�������P�M�������U�R�M������E� �j�M�-���E��j�M����E��]Ë�9�N�c�x������� ������������������������������������������������������������������������������������������̋�U��pu���@u"�pu���pu�EP�M������E���MQ�UR��������E]�����������������������̋�U����EP�M������pu��U�}� t�}�?tq�}�Xt��   �E�Pj�MQ��������E�   �pu���pu�M��4�����thTz�M������E�   ��E�Ph�{�MQ�f������E�n�pu���puj �M��h���Pj �E�P�M�Q�5�����P�M��S����U�R�EP�������E�$�M�Q�M������E��U�R�EP�������E��]����������������������������������������������������������������������������������̋�U���(�M������pu��M܃}�B��  �U���8��$�$��MQj�UR�������E�  h�{�M������M�������u
j �M�������EP�M�� ����pu���pu�M������P�U�R�EP��������E�>  �pu�Q��$t;�pu�H��u�URj�EP��������E�  �j�M�� ���E��   �pu���pu�pu��E؃}�C��   �M������$�|��pu���pu�MQ�UR�������E�   �pu���puj�MQ�UR� ������E�u�pu���puj �M��.���Pj �MQ�U�R�������P�EP�������E�9�MQj�UR�
������E�"j�M������E��EP�MQ�n������E��]ÍI f�������
� ���_������� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��� �pu��M�}�XtD�}�Zt�`�pu���pu������t	�E�H!��E��{�E�P�M�=����E��   �pu���puhTz�M�����E��   �U�R�������M����������   �pu��M�}� t�}�@t`�}�Zt�v�U�R�M�i����E�   �pu���pu������t	�E��{��E�{�M�Q�U�R�M��'���P�M�"����E�>�pu���pu�M�Q�M�����E� j�M�E����E���U�R�M������E��]��������������������������������������������������������������������������������������������̋�U���,�E�   �M������M��������  �pu���@��   �pu���Z��   �}� t	�E�    �
j,�M�������pu�����   �pu���0�M�x3�}�	-�pu���pu�E�P�M�Q�du����P�M��5����k�pu�U�M������P�E�P�Z������pu+M��~�du�n�����u�U�R�du�-����E�P�M�������pu;M�u
j�M������j�M��o����������U�R�M�>����E��]����������������������������������������������������������������������������������������̋�U���(�pu���tg�pu���Zu'�pu���pu�M������P�M�����E�^�0j)�UR�E�P������Ph�{�M�Q��������������E�,�*j)�URj�E�Ph�{�M�譻�����$����������E��]�������������������������������������������������������̋�U���x�pu����Y  �pu��E��pu���pu�E� �E������M�������U��U��E���C�E��}��  �M���h��$�<�h�|�M��p����-  h�|�M��^����  h�|�M��L����	  h�|�M��:�����  h�|�M��(�����  hx|�M�����hp|�M�������  �E����E��  �pu��U��E�E��pu���pu�U��U��}�Y�&  �E������$����E������  hh|�M������  h`|�M�������   hT|�M��v�����   hH|�M��d�����   h<|�M��R����   h0|�M��@����   h$|�M��.����   �pu���pu�E�P�l�����P�M��\����M��������t�M�Q�M������E�~  �R�UR�E�P������Ph|�MQ��������E�R  �pu���puj�M�������h|�M������QhTz�M������B�pu���pu�M�Q�������P�M�起���M��$�����t�U�R�M�X����E��  �}����   �E��E��M���C�M��}���   �U���$��$���M�Qh|�U�R�$�����P�M��B����e�E�Ph�{�M�Q������P�M��"����E�U�U��E���E�E��}�w/�M���L��$�D��E�Ph|�M�Q������P�M��۶���M�J�����u�URj �E�P�P�����P�M��ڽ���M�Q�M�c����E��   ��   �M������UR�M��B����}��uF�M������E�P�M�Q�U�R��������M�������uh8w�M��|����E�P�M������E�}�M������tA�M���t$h�{�M�������U���th�{�M��5�����E���th�{�M������M�Q�U�R�EP�������E���MQj�UR��������E��]Ë� �2�D�V�h���z�������   










	�I ������,�>�P�����b�t��� 	

��������� �I ���     ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���8�k�����t�/�����u	�E�   ��E�    �EЉE��M�������pu��U̡pu���pu�M̉Mȃ}�Y��   �U���4��$���pu���puh�|�M�ó���E�   h�|�M��:����kh�|�M��+����\h�|�M������Mh�|�M������>h�|�M�������/�����E��U�R������Ph�|�E�P������P�M��$����M������}� t�M�Q�M��
����U�R蔵����P�M������E�P�M�����E��]Ë�2�V�e�t��������� ���������������������������������������������������������������������������������������������������������������������������������̋�U��EP�y������E]����������̋�U����M������pu�����   �pu��E�M��0�M�}�wH�U��$�D�h}�M������>h }�M������/�-h�|�M�������hx|�M�������j�M�B����E�~�pu��M�pu���pu�E�E�M��1�M�}�w/�U���l��$�d��M�Qh|�U�R������P�M��ԯ���E�P�M�����E��j�M������E��]�u�u�������������� �    ��������������������������������������������������������������������������������������������̋�U����   �pu���u�URj�EP�������E�  �pu���6|�pu���9~ �pu���_tj�M������E��  �pu���6�U��pu���pu�}�)u[�pu���t2�pu���=�M��pu���pu�}�|�}�~�E�������EPj�MQ�Q������E�M  ��}� |�}�~�E������}��uj�M�#����E�   �M������UR�M������E����  �M�Qh�y�U�R������P�M��ҭ���pu���t5�U�R�E�P�M�Q�������Pj �U�R�6�����������P�M�蓭����E�Pj�M�Q������P�M��v����pu���t1�pu���@u�pu���pu�j�M�M����E�J  ��M�Qj�UR�2������E�.  �o�����t�E�P������P�M�� �����M�Q������P�M��j����U���tS�������t5�E�P�M�Q�U�R藹����Pj �E�P�H������������P�M�襬����M�Q�j�����P�M�����觱����t)�U�R��x���P�M�Q�b�����������P�M��^������p���R�A�����P�M�������M購����u.j)��`���P�M�Qj(��h���R���������&���P�M��
���j hPuj踳������\�����\��� t��\����������0����
ǅ0���    ��0����E��M�Q�U�R������j)��D���P��T���Q�s�����Pj(��L���R������������P�M�蠲���˴����t�E���t�M�Q�M�胲���\�����t��<���R������P�M��b������4���P�������P�M������}� t�M�Q�M������j�M�����E��U�R�M讽���E��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����pu�����   �pu���6|�pu���9~�pu���_uo�UR�M������M�������u$�M������u�M�-�����u�EP�M��|����M�Ź����u�MQ�M��d����U�R�EP�r������E�   �=j �MQ�UR�EP�M�Q�������U3���*��P�M�Q�UR蛬�����E�n�lj�M�������EP�M��E����M�=�����u�MQ�M��ܯ���M�%�����u"�M������u
j �M������UR�M�讯���E�P�M�7����E��]�������������������������������������������������������������������������������������������������̋�U���0�M�������pu���pu�pu��UЀ}�At�}�Bt;�}�Ctq�   �} u�E���&��ɀ�9��%�U�
�pu���pu�  �} tj�M�����E�}  �M�j>�M��>����pu���pu�N  �E� %�pu���pu�4  �pu���t�pu�Q��uj�M�5����E�  �} tj�M�����E��   �pu���0���pu�B�LЉM�pu���pu�}�v/j,�M������E�3�QP�M�����P�U�R�M������P�M�触��j>�E�P�M�����P�M�萦���pu���$u�pu���pu�j^�M�Q�M��x���P�M��\����pu���t�pu���pu�
j�M������M�������U�R�M�۸���E��M�����E��]����������������������������������������������������������������������������������������������������������������������������������������̋�U���$  �M��j����E� �pu����  �pu���$u8�MQ�U�R�EP�M�Q�P������M�覵����u�U�R�M�ڷ���E�  �pu��pu�3҃�A����+��+ʉM�M�������M�������E�   �E艅����������t������tw��������   �  �ũ����tW������tN�M��	�����u/j������P�M�Qj �U�R�M��������!���P�M��a����j�������P�M�������   �`�����tN�M�譴����u/j	������P�E�Pj �M�Q�M��(����������P�M������j	�x�����P�M������`������tN�M��T�����u/j�N�����P�U�Rj �E�P�M���������l���P�M�謣���j������P�M��@�����E�    �}� t|�pu���pu�pu���$u8�MQ�U�R�EP�M�Q�l������M��³����u�U�R�M������E�  �pu��pu�3҃�A����+��+ʉM�}� �)����pu���t�pu���pu�}���  �EP�M������M�Q�U�R�M������P�M�跢���M��&�����u)�E�P��|���Qj �U�R�M�����������P�M�肢���M�������u,�E�P��l���Qj ��t���R�M��m������o���P�M��J����E���  �} tj�M�9����E�  �M��tz�U�Rh�y��d���P�߷����P�M�������pu���t,�E�P��T���Q��\���R��������������P�M��ơ����E�Pj��L���Q������P�M�覡���%�pu���t��D���Q������P�M�� ����pu���uj�M��A����-�pu��pu���pu��@tj�M�L����E�  �R�����t[�M��������������t�B�} tj�M�����E�t  �U�R��4���P��<���Q躭�����������P�M��נ���#�U����u��,���P莭����P�M��3����M��t!�U�Rh}��$���P�k�����P�M�艠���M��t!�U�Rh}�����P�B�����P�M��`����} ��   �M�Ű������   �M������u�M詰����t:�M�������t�MQ�M�������URj �����P������P�M������@�MQ������Rj �����P�MQj �����R�^�������������������P�M��ڦ���*�M�!�����u�EPj ������Q�$�����P�M�讦���M������U���t�M��i����E�P�M�����E��   �j�M�[����E�   �   �} ux�M謯����ul�M�������u�M蔯����t�MQj�UR�������E�u�9�EP�MQj ������R�EPj������Q����������������������E�:�8�} u%�M�.�����u�URj�EP�������E��j�M�����E��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����pu����  �} t]�pu���XuO�pu���pu�M�������thTz�M荝���E��   ��URh�{�EP�*������E��   �pu���Yu%�pu���pu�MQ�UR�������E�   �EP�M�Q蚰�����M������t �U�Rh4}�E�P辱����P�M��ܛ���*�M������t�M�Qh$}�U�R蒱����P�M�谛���E�P�M�_����E���MQj�UR�������E��]��������������������������������������������������������������������������������̋�U���   �pu����s  �B����E��}� }�E�    �}� u>j]�U�Rj�E�Pj[�M��������|����������P�MQ�a������E�  �  �M������M�_�����th8w�M��ϵ���M�薪����tR�U��E����E���tB�pu���t5j]�E�Pj �M�Q�������Pj[�U�R����������_���P�M��i���뢋M谪����u^�M�������t�E�P�M�Q�M�5���P�M������7�U�R�E�Pj)�M�Q�URj(�E�P��������������������P�M��י���M�Q�U�R�2������M�������E�P�M�n����E�   �   �M������uSj]��|���Qj�U�RhD}�E�P�MQj(�U�R��������� �������������n���P�EP�������E�?�=j]��d���Qj��l���Rj[��t����[������������-���P�EP衭�����E��]��������������������������������������������������������������������������������������������������������������������������������������������������̋�U���j'�EPj �M�Q�������Pj`�U�R����������U����E��]�����������������������̋�U���j�M�����Pj �M�� ���P�EP�ӣ�����E��]���������������̋�U��j*�EP�MQ�UR�=������E]����������������̋�U��j �EP�MQ�UR�������E]����������������̋�U��j&�EP�MQ�UR�ݷ�����E]����������������̋�U��j�EP��������E]��������̋�U��j �EP�������E]��������̋�U��j �EP�������E]��������̋�U��EP�MQ诫�����E]������̋�U��Q�pu��M��}� t)�}�At�0�pu���puhH}�M跗���E�j�M�����E�j�M�����E��]���������������������������������̋�U���@�EP�M�������M��7������b  �pu����Q  �E�P�M�Qj �U�R�E�P�K�����������������P�M������M��������  �pu���@��   hT}�M������M�趥������   �pu�����   �pu���@txj'�M�Q�U�R������Pj`�E�P���������|���P�M�膜���pu���@u�pu���pu�M��<�����t�pu���@thP}�M��N����Z����M�������t �pu���u
j�M��И��j}�M��d����pu���@u�pu���pu�'�M��Ť����t�U�Rj�E�P������P�M�觔���M�Q�M�V����E��]����������������������������������������������������������������������������������������������������������������̋�U��EP�[������E]����������̋�U���j �M������Pj �M������P�EP賟�����E��]���������������̋�U����EP�M��k���hT}�M��Ӯ���M�Q辿����P�M�贚��j}�M�������pu���@u�pu���pu�U�R�M�����E��]��������������������������������̋�U���,j hPuj�ښ�����E��}� t�M������E���E�    �EԉE�M�Q�U�R蟓�����EP�M�Qj �U�R�E�P��������������������P�M�跒���M�Q�M�f����E��]������������������������������������������������̋�U�졀u�������]����������̋�U�졀u%   �����]��������̋�U�졀u�������]����������̋�U�졀u�������]����������̋�U�졀u�������]����������̋�U�졀u��`3Ƀ�`����]�������̋�U�졀u%�   �����]��������̋�U�졀u%   �����]��������̋�U�졀u%   �����]��������̋�U�졀u%   ]���������������̋�U�졀u%    ]���������������̋�U�졀u% @  ]���������������̋�U�졀u% �  �����]��������̋�U�졀u%   �����]��������̋�U��蘘����t�E���w���M���w��]���������������������̋�U�졀u�������]����������̋�U��EP�MQ�Pu�T���]�������̋�U����M�E������E�} t�MQ�U��Ѓ���   ��   �} w�E   �M�Q;U��   �}   v3��   jhPuh  �~������E��}� t�M�������E���E�    �E��E��}� tA�M�y t�U�B�M���U�E��B��M�U��Q�E�M��H�   +U�E�P�3��!��M�Q+U�E�P�M�Q�E�H�D
��]� ���������������������������������������������������������������������̋�U��Q�M��E��     �E���]�������̋�U����EP�MQ�UR�M��ڦ����輽���E��]���������������������̋�U����EP�MQ�UR�M��s������}����E��]����������������������̋�U����EP�MQ�UR�M��E������=����E��]����������������������̋�U��Q�M��E��     �M��Q�� ����E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�E���]�����������������������������������������������������̋�U��Q�M��E��H�� ����U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M��tj�UR�M��H����E���]� ������������������������������������������������������������̋�U��Q�M��E��M���I�H�E���]� �������������̋�U����M��} tdj hPuj�q������E��}� t�EP�M������E���E�    �M��U��E����Ƀ�������   �U��B% �����M��A��U��B% ����M��A�U��    �E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�E���]� ���������������������������������������������������������������������������������������̋�U��Q�M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�} t�MQ��"  ��P�UR�M������E���]� �������������������������������������������������������������������̋�U���V�M�E�H�� ����U�J�E�H�������U�J�E�H�������U�J�E�H�������U�J�E�H�������U�J�E��     �M�Q�������E�P�M�Q�������E�P�M�Q�������E�P�M�Q������E�P�M�9 ��  �U������  �E�    �U��E���M����E��M�����  �M���M;���   �U����_��   �U����$��   �U����<��   �U����>��   �U����-tw�U����a|�U����z~]�U����A|�U����Z~C�U����0|�U����9~)�U�����   |�U�����   ~	者����t�U����U���E�H�� ������U�J�   ������E�P�M�Q�M������U����t<�U�E���M�	���u�;�t�U�B% ������M�A�U��    �!�M�躷����u�E�H�� ������U�J��E�H�� ������U�J��E�H�� ������U�J�E�^��]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�졀u%   ]���������������̋�U���$�XD3ŉE��M܍E��E��M܋Q�� ����E܉P�M��    �U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%����M܉A�U�� �E����E�j j
�MQ�UR蹪����0�� �M��j j
�UR�EP�,����E�U�MMu��U��E�+й   +�Q�U�R�M��~����E܋M�3�������]� ����������������������������������������������������������������������������������������̋�U���(�XD3ŉE��M؍E��E܋M؋Q�� ����E؉P�M��    �U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%����M؉A�U�� �E� �} |�} s�E��E�؋M�� �ىE�M�U܃��U�j j
�EP�MQ� �����0�� �U܈j j
�EP�MQ�s����E�U�UUu��E��t�M܃��M܋U��-�E܍M�+��   +�R�E�P�M������E؋M�3��<�����]� ��������������������������������������������������������������������������������������������������������̋�U����M��E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�}t�}t	�E�    ��E�E��M����   �U��B% �����M��A�U��    �}u.�EP�������M���U��: u�E��H�� ������U��J�E���]� �����������������������������������������������������������������������̋�U��Q�M��E��H����3�������]���������������̋�U��Q�M��E�3Ƀ8 ������]������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H��   �U��J�E���]��������������̋�U��Q�M��E��@������]�������̋�U����M��M��x�����u�E��H��	��t	�E�   ��E�    �E���]��������������������̋�U��Q�M��M��*�����u�E��H��   �U��J��]���������������������̋�U����M��M�������u�E��H��
��t	�E�   ��E�    �E���]��������������������̋�U��Q�M��E��H��   �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H��   �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H��    �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H�� @  �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H�� �  �U��J��]�����������������̋�U��Q�M��M��
�����t3���E���U����ȋ�Ћ�]�����������������̋�U��Q�M��M��ʍ����t2���E���U����ȋB�Ћ�]����������������̋�U����M�M�舍����uX�} u*�M��۠�����Ej hPu�EP襄�����E��M��M�} t �U�E�L�Q�UR�M��ȗ���E��E��  ��} t�M� �E��]� �������������������������������������������̋�U��Q�M��M��ڌ����t�E��EP�MQ�U���M��	��B�Ћ�]� ����������������������̋�U����M�E�P�M��Ȏ���MQ�M��w����U�R�M诎���E��]� ����������������������̋�U����M�E�P�M��x����MQ�M������U�R�M�`����E��]� �����������������������̋�U����M�E�P�M��(����MQ�M�臂���U�R�M�����E��]� �����������������������̋�U����M�E�P�M��؍���MQ�M������U�R�M������E��]� �����������������������̋�U����M�E�P�M�舍���MQ�M��~���U�R�M�p����E��]� �����������������������̋�U����M��} t_j hPuj�1������E��}� t�EP�M��R�M��O����E���E�    �E��M��U��: u�E��H�� ������U��J��E��H�� ������U��J��]� ������������������������������������̋�U����M��M��Љ����tb�E��tZ�M��4�����t�MQ�M��m����?j hPuj�X������E��}� t�UR�M�螕���E���E�    �E�P�M��S����E���]� ���������������������������������������������̋�U����M��M�� �����tu�} to�E���te�M��|�����t�UR�M�螱���Kj hPuj血�����E��}� t�EP�  ��P�MQ�M������E���E�    �U�R�M�萐���E���]� ������������������������������������������̋�U��Q�M��M��b�����tG�M�Έ����t�M�8���P�M��|���(�M�诈����t�EP�M��(x����M�R�M�� ����E���]� ��������������������������̋�U����M��M����������   �} ��   �M��>�����t�EP�M������j�M蚨����t�M莨����u@j hPuj�J�����E��}� t�MQ�M������E���E�    �U�R�M��F�����M�A���P�M��${���E���]� ���������������������������������������������̋�U��Q�M��M�������tC�M��n�����u�}t�}u�EP�M��դ����} u��MQ荘����P�M�褎���E���]� ������������������������������̋�U����M��M��n�����t3�M�s�����u'�M�U����E��E�%�   �M��Q�� ���ЋE��P�E���]� ���������������������������̋�U��Q�M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M��tj�UR�M��X����E���]� ������������������������������������������������������������̋�U��Q�M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�MQ�  ��P�UR�M��E����E���]� ���������������������������������������������������������̋�U��Q�M��E��M���I�H�E���]� �������������̋�U����M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�} tXj hPuj��z�����E��}� t�MQ�M��\����E���E�    �U��E��M��9 u�U��B% ������M��A��U��B% ������M��A�E���]� ������������������������������������������������������������������������������̋�U��Q�M��E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�E%�   �M��Q�� ���ЋE��P�}u0�MQ�U������U���E��8 u�M��Q�� ������E��P�	�M��    �E���]� ������������������������������������������������������������������̋�U����M�E�8 tj�M������  �} ��   �} ��   �M�M��}� t�}�t�u�U�B% ������M�A�   j hPuj�_x�����E��}� t�U�P�M�裌���E���E�    �M�U��E�8 u�M�Q�� ������E�P�[j hPuj�x�����E��}� t�MQ�UR�M��V����E���E�    �E�M��U�: u�E�H�� ������U�J��E�H�� ������U�J��]� ����������������������������������������������������������������������������������������̋�U��Q�M��E�3Ƀ8	������]������̋�U��Q�M��E�� �����E���]�������̋�U����M�M���r����uf�M�����uZj hPuj��v�����E��}� t�EP�M�趁���E���E�    �M��M��}� t�U����M��U��M�U��T��E��]� �����������������������������������������̋�U��Q�M��} |�}	~j�M耮���E�;�9�E��8�t
�M��U;~j�M�]����E���E�M��T�R�M�����E��]� ��������������������������̋�U��Q�M��E�� \}�E���]�������̋�U��Q�M��M�趋���E�� l}�M��U�Q�E���]� �������������������̋�U��Q�M��   ��]��������������̋�U��Q�M��E��@��]�������������̋�U��Q�M��E;Es�M�U��B��M���M�E��]� �����������������̋�U����M��M������E�� |}�} tP�} tJj hPu�MQ�t�����E��U��E��B�M��U�Q�E��x t�MQ�UR�E��HQ�S  ����U��B    �E��@    �E���]� ������������������������������������������������̋�U��Q�M��E��@��]�������������̋�U����M��E��x t�M��Q�E��H�T
��U���E� �E���]����������������������������̋�U��Q�M��E��HQ�U��BP�MQ�UR�n�������]� ������������������̋�U��Q�E+E�E��M;M�~�U��U�EP�MQ�UR�"  ���EE��]���������������������̋�U����M��M��4����E�� �}�} t#�M�7�����t�M�*�����u	�E�    ��M�M��U��E��B�E���]� ����������������������������������̋�U����M��E��x t�M��I豎���E���E�    �E���]��������������̋�U����M��E��x t�M��I蚈���E���E� �E���]�����������������̋�U����M��E��x t�MQ�UR�E��H�U����E���M�M��E���]� ��������������������̋�U��Q�M��M������E�� �}�M��U�Q�E��H����Ƀ�����U��J�E���]� ��������������������������̋�U��Q�M��E��@��]�������������̋�U��Q�M��E��x��,"�}��]�����������������̋�U��Q�M��E��xujh�}�MQ�UR�܏������E��]� ���������������������������̋�U��j�h��d�    P�XD3�P�E�d�    �4v��uM�4v���4v�E�    j ��u薗��j�v芗��j�v�~���j�v�r����E������} |�}}�Ek��u��v�M�d�    Y��]��������������������������������������������������������̋�U��Q�M��M������E�� �}�M��U�Q�E��M�H�U��B�����E���]� ����������������̋�U��QV�M��E��x }.�M��Q�E��H���Ћ��M��Q�E��H������M��q�U��B^��]��������������������̋�U����M��E��H�U��B��ȋB�ЈE��M���u�U��B�M��I��B�ЈE��E���]������������������������̋�U����M��EP�MQ�U��B�M��I��B�ЉE��M�;Ms�UR�E�P�M��Q�E��H��B�����E���]� ����������������������̋�U��Q�E�    �	�E���E�M���t�E����E���E���]����������������������������̋�U��Q�E�    �	�E����E��M�;Ms�UU��EE���
�݋�]��������������������������̋�U��} u3��G�E���Et.�M���t$�E��U�;�u�M���M�U���U�ǋE� �M�+�]�������������������������SVW�T$�D$�L$URPQQh�d�5    �XD3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�!����   �C�+n���d�    ��_^[ËL$�A   �   t3�D$�H3�蝏��U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�~��3�3�3�3�3���U��SVWj j hwQ蕡��_^[]�U�l$RQ�t$������]� ��������������������������������������������������������������������������������������������̋�U��E�8v]�����������������̋�U��j�hX.h"�d�    P���SVW�XD1E�3�P�E�d�    �e��E�    �EP�MQ����E��E������;�U���M��U�3���  ���Ëe�}�  �uj� ��E�    �E������E�M�d�    Y_^[��]������������������������������������������̋�U���L�E�    �} t�} u3��(  �} t�} v3��Mf�3҃} �U�}� uhp~j jEh�}j��i������u̃}� u.�P����    j jEh�}h�}hp~�}��������  �MQ�M��s���} �  �M���h����z uj�E�;EsG�MM�f��Ef��MM����u�E��E؍M�蠈���E��O  �M����M��U���U뱋E��EԍM��v����E��%  �  �MQ�URj��EPj	�M��]h����QR�ܒ�E��}� t�E����EЍM��+����E���  �����zt*�A���� *   3ɋUf�
�E������M�������E��  �E�E��M�M��	�U���U�E��M����M���tk�U����ta�M���g��P�M��R��i������t@�E��H��u,迆��� *   3ҋEf��E������M��t����E��#  �	�M���M��|����U�+U�U܋EP�MQ�U�R�EPj�M��Eg����QR�ܒ�E��}� u*�M���� *   3��Mf��E������M������E��   �U��U��M������E��   �   �M���f��� �x u�MQ�'������E��M�踆���E��j�`j j j��URj	�M��f��� �HQ�ܒ�E��}� u!豅��� *   �E������M��n����E�� ��U����U��M��V����E���M��I�����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EP�MQ�UR�EP�ޕ����]�����������������̋�U��=u uh�W�EP�MQ�UR�و������j �EP�MQ�UR迈����]�����������������������������̋�U���L�E�    �} u�} t�} t�} w	�E�    ��E�   �EĉE��}� u!hj h�   h�}j�e������u̃}� u3蒃���    j h�   h�}h�~h��x�����   ��  �} tY3ҋEf��}�tK�}���tB�}v<�M��9�Hs��H�U��	�E���E��M���Qh�   �U��R�k������} t	�E�     �MQ�M��^n���U;Uv�E�E���M�M��U��U�����;E�Ƀ��M�u!h�~j h  h�}j�d������u̃}� u@萂���    j h  h�}h�~h�~��w�����E�   �M��/����E���  �M��+c��P�E�P�MQ�UR袓�����E�}��ux�} tX3��Mf��}�tJ�}���tA�}v;�U��9�Hs
��H�E��	�M���M��U���Rh�   �E��P�7������́����MЍM�葂���E��/  �U���U�} ��   �E�;E��   �}���   3ɋUf�
�}�tK�}���tB�}v<�E��9�Hs��H�M��	�U���U��E���Ph�   �M��Q蛌�����U�9U����E�u!h�~j h  h�}j�wb������u̃}� u=������ "   j h  h�}h�~h�~�Lv�����E�"   �M�蘁���E��9�U�U��E�P   3��M�Uf�DJ��} t�E�M��U��UȍM��]����Eȋ�]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�5�����]�����������̋�U���4�} t�} v	�E�   ��E�    �E�E�}� uh��j jh��j�`������u̃}� u0����    j jh��hp�h���nt�����   �K  �} ��   �U� �}�tI�}���t@�}v:�E��9�Hs��H�M��	�U���U��E�Ph�   �M��Q������3҃} �U��}� uhЗj jh��j��_������u̃}� u0�S~���    j jh��hp�hЗ�s�����   �  �M�M��U�U��}� v�E����t�U����U��E����E��܃}� ��   �M� �}�tH�}���t?�}v9�U��9�Hs
��H�E��	�M���M܋U�Rh�   �E��P� ������(���t3�t	�E�   ��E�    �E؉E�}� uh�j j h��j��^������u̃}� u0�H}���    j j h��hp�h��r�����   �{  �U��E��
�U���M����M��U���U��t�E����E�t�̓}� ��   �M� �}�tH�}���t?�}v9�U��9�Hs
��H�E��	�M���MԋU�Rh�   �E��P�����������t3�t	�E�   ��E�    �EЉE�}� uhX�j j*h��j�]������u̃}� u-�:|��� "   j j*h��hp�hX��q�����"   �p�}�th�}���t_�U+U���;UsQ�E+E����M+�9�Hs��H�U���E+E����M+ȉM̋U�Rh�   �E+E��M�TR�
�����3���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���8�E؉E�3Ƀ} ���Mԃ}� uhmj jph�lj��[������u̃}� u.�Xz���    j jph�lhX�hm�o��������P  �} t�} u	�E�    ��E�   �ẺEЃ}� uh�j jsh�lj�\[������u̃}� u.��y���    j jsh�lhX�h��4o���������   �}���v�U��B����	�E��M�H�U��BB   �E��M�H�U��E��MQ�UR�EP�M�Q�U���E��} u�E��y�}� |V�U��B���M��A�U��z |"�E��� 3ҁ��   �UȋE�����U��
��E�Pj �&o�����Eȃ}��t�E���MM�A� �U��z }�����������]��������������������������������������������������������������������������������������������������������������������������̋�U����EPj �MQ�UR�EPh[�������E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQh[��8�����E��}� }	�E�������U��U��E���]������������������������̋�U��� �E�����3��} ���E��}� u!h8�j h�   h�lj��X������u̃}� u1�Tw���    j h�   h�lh�h8��l���������  �} t�} v	�E�   ��E�    �U�U�}� u!h��j h�   h�lj�RX������u̃}� u1��v���    j h�   h�lh�h���'l��������d  �MQ�UR�EP�MQ�URh����}�����E��}� }U�E�  �}�tI�}���t@�}v:�M��9�Hs��H�U��	�E���E�M�Qh�   �U��R菁�����}��uu3�t	�E�   ��E�    �M�M��}� u!h��j h�   h�lj�UW������u̃}� u.��u��� "   j h�   h�lh�h���*k��������j�}� |a�}�t[�}���tR�E���;EsG�M����U+�9�Hs
��H�E���M����U+щU��E�Ph�   �M��U�D
P譀�����E���]���������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP��n����]���������������̋�U���,�E������E�    3��} ���E�}� u!h8�j h  h�lj�U������u̃}� u1�t���    j h  h�lh\�h8��pi��������  �} u�} u�} u3���  �} t�} v	�E�   ��E�    �U�U��}� u!h��j h  h�lj�U������u̃}� u1�s���    j h  h�lh\�h����h��������|  �M;M��   �Gs����U��EP�MQ�UR�E��P�MQh���~z�����E��}��u~�}�t\�}���tS�U��;UsH�E���M+�9�Hs��H�U���E���M+ȉM�U�Rh�   �E�M�TR�~�����r���8"u
�r���M������  �`�r����U��EP�MQ�UR�EP�MQh����y�����E��UU�B� �}��u"�}�u�Lr���8"u
�Br���M������Y  �}� ��   �U� �}�tI�}���t@�}v:�E��9�Hs��H�M��	�U���U��E�Ph�   �M��Q�<}�����}��uu3�t	�E�   ��E�    �E܉E�}� u!h��j hB  h�lj�S������u̃}� u.�q��� "   j hB  h�lh\�h����f������������z�}�t\�}���tS�U���;UsH�E����M+�9�Hs��H�U���E����M+ȉM؋U�Rh�   �E��M�TR�Z|�����}� }	�E�������E��EԋEԋ�]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�MQ��H����]�����������̋�U����EPj �MQ�UR�EPh����v�����E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQh���v�����E��}� }	�E�������U��U��E���]������������������������̋�U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP�@   �E��j �MQ�UR�EP�MQ�$   �E��E���]��������������������������̋�U���03��} ���E�}� uht�j jfh��j��O������u̃}� u0�Nn���    j jfh��h��ht��c�����   ��  3�;U��؉E�uhX�j jgh��j�jO������u̃}� u0��m���    j jgh��h��hX��Bc�����   �  �U� �}�tI�}���t@�}v:�E��9�Hs��H�M��	�U���UԋE�Ph�   �M��Q��x����3҃} ��;U��؉E�uh��j jih��j�N������u̃}� u0�+m��� "   j jih��h��h���b�����"   ��  �}r�}$w	�E�   ��E�    �UЉU܃}� uh��j jjh��j�-N������u̃}� u0�l���    j jjh��h��h���b�����   �O  �E�    �M�M��} t �U��-�E����E��M����M��U�ډU�E��E�E3��u�U�E3��u�E�}�	v�M��W�U��
�E����E���M��0�U��
�E����E��M����M��} v�U�;Ur��E�;Erl�M� �U�;U��؉E�u!h��j h�   h��j�#M������u̃}� u0�k��� "   j h�   h��h��h����`�����"   �E�U�� �E����E��M���U�E��M���E�M��U����U��E���E�M�;M�r�3���]� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�}
u�} }	�E�   ��E�    �E�P�MQ�UR�EP�MQ������]�����������������̋�U��j �EP�MQ�UR�EP�T���]������������������̋�U��Q�}
u�} |�} s	�E�   ��E�    �E�P�MQ�UR�EP�U�M�   ��]�����������������������̋�U���8�UЉM�3��}� ���E�}� u!ht�j h>  h��j�J������u̃}� u3�%i���    j h>  h��h �ht��x^�����   �,  3�;U���؉E�u!hX�j h?  h��j�;J������u̃}� u3�h���    j h?  h��h �hX��^�����   ��  �U�� �}��tI�}����t@�}�v:�EЃ�9�Hs��H�M��	�UЃ��ŰE�Ph�   �Mԃ�Q�s����3҃} ��;U���؉E�u!h��j hA  h��j�tI������u̃}� u3��g��� "   j hA  h��h �h���I]�����"   ��  �}r�}$w	�E�   ��E�    �UȉU܃}� u!h��j hB  h��j��H������u̃}� u3�tg���    j hB  h��h �h����\�����   �{  �E�    �MԉM��} t+�U��-�E����E��M����M��U�ڋE�� �؉U�E�M��M�U3�PR�MQ�UR�4g���E�E3�QP�UR�EP�d���E�U�}�	v�M��W�U��
�E����E���M��0�U��
�E����E��M����M��} w�} v�U�;U�r��E�;E�rl�M�� �U�;U���؉E�u!h��j hf  h��j�G������u̃}� u0�;f��� "   j hf  h��h �h���[�����"   �E�U�� �E����E��M���U�E��M���E�M��U����U��E���E�M�;M�r�3���]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�U�M�B���]����������������̋�U���l�XD3ŉE��E�    �E�    �} t�} u3��H  3��} ���EЃ}� uh��j jfhH�j�E������u̃}� u.�3d���    j jfhH�h�h���Y���������  �UR�M��rO���} �.  �M���D��� �x ��   �M�;Msp�U�=�   ~"��c��� *   �E������M��d���E��  �MM��U���M��E���E��u�M��MȍM��Md���E��M  �U����U�눋E��EčM��,d���E��,  �  �M��#D������   ��   �} v�UR�EP�2  ���E�M�Qj �UR�EP�MQ�URj �M���C��� �HQ�ؒ�E��}� t3�}� u-�UU��B���u	�M����M��U��U��M��c���E��  �b��� *   �E������M��mc���E��m  ��  �E�Pj �MQ�URj��EPj �M��NC����QR�ؒ�E��}� t�}� u�E����E��M��c���E��  �}� u�����zt"�&b��� *   �E������M���b���E���  �M�;M�  �U�Rj �M���B��� ���   Q�U�Rj�EPj �M��B����QR�ؒ�E�}� t�}� t"�a��� *   �E������M��ob���E��o  �}� |�}�v"�a��� *   �E������M��Ab���E��A  �E�E�;Ev�M��M��M�� b���E��   �E�    ��U����U��E����E��M�;M�}4�UU��E��LԈ
�UU����u�M��M��M���a���E���   벋U���U������E��E��M��a���E��   �   �M��A����y u�UR�cn�����E��M��qa���E��t�j�E�Pj j j j��MQj �M��\A����BP�ؒ�E��}� t�}� t�^`��� *   �E������M��a���E���M����M��M��a���E���M���`���M�3��e����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E���E��M�M��U����U�t�E����t�U����U����}� t�E����u�E�+E������E��]�������������������������������������̋�U��EP�MQ�UR�EP�^W����]�����������������̋�U��j �EP�MQ�UR�0W����]�������������������̋�U���,�E�    �} t�} w�} u�} t	�E�    ��E�   �E�E��}� u!h8�j h3  hH�j� ?������u̃}� u3�]���    j h3  hH�h�h8���R�����   �  �} tU�U� �}�tI�}���t@�}v:�E��9�Hs��H�M��	�U���U��E�Ph�   �M��Q�h�����} t	�U�    �E;Ev�M�M���U�U܋E܉E�����;M�҃��U�u!h�~j h?  hH�j�.>������u̃}� u3�\���    j h?  hH�h�h�~�R�����   �  �MQ�U�R�EP�MQ�tU�����E�}��ug�} tU�U� �}�tI�}���t@�}v:�E��9�Hs��H�M��	�U���U؋E�Ph�   �M��Q�lg�����\��� �  �U���U�} ��   �E�;E��   �}���   �M� �}�tH�}���t?�}v9�U��9�Hs
��H�E��	�M���MԋU�Rh�   �E��P��f�����M9M���ډU�u!h��j hW  hH�j��<������u̃}� u0�B[��� "   j hW  hH�h�h���P�����"   �(�M�M��E�P   �UU��B� �} t�E�M��E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ��d����]�����������̋�U���4�} t�} v	�E�   ��E�    �E�E�}� uhx�j jh��j�;������u̃}� u0�Y���    j jh��h��hx���N�����   �\  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9�Hs��H�U��	�E���E��M���Qh�   �U��R�pd����3��} ���E��}� uhЗj jh��j�M:������u̃}� u0��X���    j jh��h��hЗ�%N�����   �  �U�U��E�E��}� v�M����t�E����E��M����M��܃}� ��   3ҋEf��}�tK�}���tB�}v<�M��9�Hs��H�U��	�E���E܋M���Qh�   �U��R�wc�����(���t3�t	�E�   ��E�    �U؉U�}� uh�j j h��j�=9������u̃}� u0�W���    j j h��h��h��M�����   �  �M��Uf�f��M���E����E��M���M��t�U����U�t�˃}� ��   3��Mf��}�tJ�}���tA�}v;�U��9�Hs
��H�E��	�M���MԋU���Rh�   �E��P�cb���������t3�t	�E�   ��E�    �EЉE�}� uhX�j j*h��j�)8������u̃}� u-�V��� "   j j*h��h��hX��L�����"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9�Hs��H�U���E+E����M+ȉM̋U���Rh�   �E+E��M�TAR�ya����3���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���<�E؉E�3Ƀ} ���Mԃ}� u!hmj h�   h(�j�C6������u̃}� u1��T���    j h�   h(�h��hm�J��������  �} t�} u	�E�    ��E�   �ẺEЃ}� u!h�j h�   h(�j��5������u̃}� u1�ET���    j h�   h(�h��h��I��������3  �U��BB   �E��M�H�U��E��}���?v�M��A�����U��E��P�MQ�UR�EP�M�Q�U���E��} u�E���   �}� ��   �U��B���M��A�U��z |"�E��� 3ҁ��   �UȋE�����U��
��E�Pj �I�����Eȃ}��tV�M��Q���E��P�M��y |"�U���  3Ɂ��   �MċU�����M����U�Rj �0I�����Eă}��t�E�� 3��M�Uf�DJ��E��x }�����������]�������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EPj �MQ�UR�EPh���?h�����E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQh����g�����E��}� }	�E�������U��U��E���]������������������������̋�U��� �E�����3��} ���E��}� u!h8�j h  h(�j��2������u̃}� u1�DQ���    j h  h(�h�h8��F���������  �} t�} v	�E�   ��E�    �U�U�}� u!h��j h  h(�j�B2������u̃}� u1��P���    j h  h(�h�h���F��������j  �MQ�UR�EP�MQ�URh��f�����E��}� }X3��Mf��}�tJ�}���tA�}v;�U��9�Hs
��H�E��	�M���M�U���Rh�   �E��P�|[�����}��uu3�t	�E�   ��E�    �U�U��}� u!h��j h  h(�j�B1������u̃}� u.��O��� "   j h  h(�h�h���E��������m�}� |d�}�t^�}���tU�M���;MsJ�U����E+�9�Hs��H�M���U����E+E��M���Qh�   �U��E�LPQ�Z�����E���]���������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP��7����]���������������̋�U���,�E������E�    3��} ���E�}� u!h8�j h9  h(�j�/������u̃}� u1�N���    j h9  h(�h�h8��`C��������&  �} u�} u�} u3��  �} t�} v	�E�   ��E�    �U�U��}� u!h��j h?  h(�j��.������u̃}� u1�tM���    j h?  h(�h�h����B��������  �M;M��   �7M����U��EP�MQ�UR�E��P�MQh��#c�����E��}����   �}�t^�}���tU�U��;UsJ�E���M+�9�Hs��H�U���E���M+ȉM�U���Rh�   �E�M�TAR�X�����L���8"u
�L���M�������  �c�zL����U��EP�MQ�UR�EP�MQh��ib�����E�3ҋE�Mf�TA��}��u"�}�u�3L���8"u
�)L���U������a  �}� ��   3��Mf��}�tJ�}���tA�}v;�U��9�Hs
��H�E��	�M���M��U���Rh�   �E��P� W�����}��ux3�t	�E�   ��E�    �U܉U�}� u!h��j hf  h(�j��,������u̃}� u1�hK��� "   j hf  h(�h�h���@��������   ����|�}�t^�}���tU�M���;MsJ�U����E+�9�Hs��H�M���U����E+E؋M���Qh�   �U��E�LPQ�9V�����}� }	�E�������U��UԋEԋ�]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�MQ�6����]�����������̋�U����EPj �MQ�UR�EPhw��_�����E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQhw��_�����E��}� }	�E�������U��U��E���]������������������������̋�U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP�@   �E��j �MQ�UR�EP�MQ�$   �E��E���]��������������������������̋�U���03��} ���E�}� uht�j jfh��j�)������u̃}� u0�H���    j jfh��h@�ht��t=�����   �  3�;U��؉E�uhX�j jgh��j�:)������u̃}� u0�G���    j jgh��h@�hX��=�����   �  3ҋEf��}�tK�}���tB�}v<�M��9�Hs��H�U��	�E���EԋM���Qh�   �U��R�R����3��} ����;E��ىM�uh��j jih��j�u(������u̃}� u0��F��� "   j jih��h@�h���M<�����"   ��  �}r�}$w	�E�   ��E�    �EЉE܃}� uh��j jjh��j��'������u̃}� u0�{F���    j jjh��h@�h����;�����   �`  �E�    �U�U��} t%�-   �M�f��U����U��E����E��M�ىM�U��U�E3��u�U�E3��u�E�}�	v�E��W�M�f��U����U���E��0�M�f��U����U��E����E��} v�M�;Mr��U�;Urn3��Mf��U�;U��؉E�u!h��j h�   h��j��&������u̃}� u0�hE��� "   j h�   h��h@�h���:�����"   �M3ҋE�f��M����M��U�f�f�E��M��U�f�f��M�f�U�f��E����E��M���M�U�;U�r�3���]� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�}
u�} }	�E�   ��E�    �E�P�MQ�UR�EP�MQ�e�����]�����������������̋�U��j �EP�MQ�UR�EP�4���]������������������̋�U��Q�}
u�} |�} s	�E�   ��E�    �E�P�MQ�UR�EP�U�M�   ��]�����������������������̋�U���8�UЉM�3��}� ���E�}� u!ht�j h>  h��j�S$������u̃}� u3��B���    j h>  h��hP�ht��(8�����   �A  3�;U���؉E�u!hX�j h?  h��j��#������u̃}� u3�mB���    j h?  h��hP�hX���7�����   ��  3ҋE�f��}��tK�}����tB�}�v<�MЃ�9�Hs��H�U��	�EЃ��E̋M���Qh�   �Uԃ�R�LM����3��} ����;E���ىM�u!h��j hA  h��j� #������u̃}� u3�A��� "   j hA  h��hP�h����6�����"   �  �}r�}$w	�E�   ��E�    �EȉE܃}� u!h��j hB  h��j�"������u̃}� u3� A���    j hB  h��hP�h���s6�����   �  �E�    �UԉU��} t0�-   �M�f��U����U��E����E��M�ًU�� �ډM�U�E��E�M3�RQ�EP�MQ��@���E�U3�PR�MQ�UR�S>���E�U�}�	v�E��W�M�f��U����U���E��0�M�f��U����U��E����E��} w�} v�M�;M�r��U�;U�rn3��M�f��U�;U���؉E�u!h��j hf  h��j�\!������u̃}� u0��?��� "   j hf  h��hP�h���15�����"   �M3ҋE�f��M����M��U�f�f�E��M��U�f�f��M�f�U�f��E����E��M���M�U�;U�r�3���]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�U�M�"���]����������������̋�U����E�E��M����MZ  t3��;�E��M�H<�M�U�:PE  t3�� �E���E��M����  t3���   ��]���������������������������������̋�U����E�MH<�M��E�    �U��B�M��T�U���E����E��M��(�M�U��B9E�s#�M�U;Qr�E�H�U�J9Ms�E���3���]�������������������������������������������̋�U��j�hx.h"�d�    P���SVW�XD1E�3�P�E�d�    �e��E�   �E�    �E�P�SO������u�E�    �E������E��   �M+M�M܋U�R�E�P�PL�����E��}� u�E�    �E������E��b�M��Q$��   ���҃��U��E������E��@�E������7�E���U؋E�3�=  �����Ëe��E�    �E������E���E������M�d�    Y_^[��]������������������������������������������������������������������������������̋�U��E�<v]�����������������̋�U���$V�<vP�/�����E�3Ƀ} ���M��}� uh|�j jDh�j�������u̃}� u0�<;���    j jDh�h�h|��0�����   �  �E�     �}� �a  h,m���E�}� ut3�t	�E�   ��E�    �U��U�}� uh��j jPh�j�������u̃}� u0�:���    j jPh�h�h����/�����   ��   hh��M�Q���E��}� ��   3�t	�E�   ��E�    �E܉E�}� uh��j jVh�j�������u̃}� uD���P� N������� :���0j jVh�h�h���Z/�������P��M�����X�U�R�R�����E���J���E��E�Ph<v�d�;E�t
�M�Q���j�UR�U���u�9���    �9��� �3�^��]����������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  �XD3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M�� $���E�    3Ƀ} �������������� u!h�nj h  h�Ej�������u̃����� uF�>8���    j h  h�Eh��h�n�-����ǅD��������M���8����D����  3��} �������������� u!hmj h  h�Ej�7������u̃����� uF�7���    j h  h�Eh��hm�	-����ǅ@��������M��R8����@����  ǅ����    �E�    ǅ����    �E�    �E�    �Uf�f�������������U���U����  ������ ��  �������� |%��������x���������D����4����
ǅ4���    ��4�����������������������ШD����������������0�����0����(  ��0����$�\~�E�   ������Q�UR������P�`  ����  �E�    �MԉM؋U؉U�E�E��E�    �E������E�    ��  ��������,�����,����� ��,�����,���wL��,������~�$�|~�U����U��-�E����E��"�M����M���U��ʀ   �U��	�E����E��K  ��������*u(�UR�1�����E�}� }�E����E��M��ىM���U�k�
�������LЉM���  �E�    ��  ��������*u�EP�Q1�����EЃ}� }�E�������M�k�
�������DЉE��  ��������(�����(�����I��(�����(���.�  ��(������~�$��~�U���lu�M���M�U���   �U��	�E����E���   �M���6u%�E�H��4u�U���U�E� �  �E��   �M���3u"�E�H��2u�U���U�E�%����E��S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    �w�����M��� �M���U���   �U��t
  ��������$�����$�����A��$�����$���7�P  ��$�����(�$��~�M���0  u	�U��� �U��E�   �EP�/����f�������M��� tW���������   ������ƅ���� �M��2��P�M��)��� ���   Q������R������P�U0������}�E�   �f������f�������������U��E�   �  �EP��.���������������� t�������y u��N�U��E�P��@�����E��P�M���   t&�������B�E���������+����E��E�   ��E�    �������B�E���������U���  �E�%0  u	�M��� �M��}��uǅ �������	�UЉ� ����� ����������MQ�".�����E��U��� ��   �}� u��N�E��M��������E�    �	�U܃��U܋E�;�����}L���������t?�M����P�������Q�������t������������������������������d�}� u	��N�M��E�   �U�����������������������������t���������t���������������ɋ�����+U����U��  �EP�-�����������eI������   3�tǅ���   �
ǅ���    �������|�����|��� u!hPEj h�  h�Ej�*������u̃�|��� uF�0���    j h�  h�Eh��hPE��%����ǅ<��������M��E1����<����  ��  �M��� t������f������f����������������E�   �  �E�   �������� f�������M���@�M��������U��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}У   ~Ah�  hEj�MЁ�]  Q��
�����E��}� t�U��U��E�]  �E���EУ   �M���M�U�B��J���p�����t����M��2��P�U�R�E�P������Q�U�R�E�P��p���Q�TIR�>#�����Ѓ��E�%�   t'�}� u!�M�����P�M�Q�`IR�#�����Ѓ���������gu+�M���   u �M����P�U�R�\IP��"�����Ѓ��M����-u�E�   �E��M����M��U�R��<�����E��  �E���@�E��E�
   �u�E�
   �l�E�   ǅ����   �
ǅ����'   �E�   �M���   t�0   f�U싅������Qf�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�?������`�����d����   �U���   t�EP�?������`�����d����   �M��� tB�U���@t�EP�)��������`�����d�����MQ�y)���������`�����d����=�U���@t�EP�S)�������`�����d�����MQ�8)����3҉�`�����d����E���@t@��d��� 7|	��`��� s,��`����ً�d����� �ډ�X�����\����E�   �E����`�����X�����d�����\����E�% �  u&�M���   u��X�����\����� ��X�����\����}� }	�E�   ��M�����M��}�   ~�E�   ��X����\���u�E�    �������E��MЋUЃ��UЅ���X����\���t{�E��RP��\���Q��X���R�a,����0��l����E��RP��\���P��X���Q��)����X�����\�����l���9~��l����������l����E���l�����U����U��g���������+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@tN�E�%   t�-   f�M��E�   �2�U���t�+   f�E��E�   ��M���t�    f�U��E�   �E�+E�+E䉅T����M���u������R�EP��T���Qj �O  ��������R�EP�M�Q�U�R�  ���E���t$�M���u������R�EP��T���Qj0�  ���}� ��   �}� ��   �U���P����E܉�L�����L�����L�������L�����~}�M��-��P�M��$��� ���   Q��P���R������P�P'������H�����H��� ǅ���������2������Q�UR������P��  ����P����H�����P����j����������R�EP�M�Q�U�R�  �������� |$�E���t������Q�UR��T���Pj �  ���}� tj�M�Q�w�����E�    �$�����������8����M��.*����8����M�3��8.����]ÍI q8qkq�q.r:r}r�s�q�q�q�q�q�q �I �r�s�r�s�s �rw�s;u>y�t�w	ty{v�y7yNu.yJy1|   	
���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�H��@t�U�z u�E����U�
�4�EP�MQ������Ё���  u�E� ������M����E�]����������������������������������̋�U��E�M���M��~!�UR�EP�MQ�Y������U�:�u���]������������������������̋�U��Q�E�H��@t�U�z u�E�M�U�
�b�E�M���M��~R�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u ��"���8*u�EP�MQj?��������랋�]�������������������������������������������������̋�U���8�E؉E�3Ƀ} ���Mԃ}� u!hmj h�   h(�j�������u̃}� u1�5"���    j h�   h(�ḧhm���������P  3��} ���EЃ}� u!h\lj h�   h(�j�I������u̃}� u1��!���    j h�   h(�ḧh\l����������   �U��BB   �E��M�H�U��E��M��A����UR�EP�MQ�U�R�_"�����E��} u�E��   �E��H���U��J�E��x |!�M��� 3�%�   �E̋M�����E����M�Qj �&�����E̋U��B���M��A�U��z |"�E��� 3ҁ��   �UȋE�����U��
��E�Pj �������EȋE���]��������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�����]�������������������̋�U��EP�MQ�UR�EP�\����]�����������������̋�U���,�E؉E�3Ƀ} ���Mԃ}� u!hmj h�  h(�j�������u̃}� u.����    j h�  h(�h�hm����������C�E��@����M��AB   �U��B    �E��     �MQ�UR�EP�M�Q�U���E��E���]����������������������������������������������������̋�U��EPj �MQh�������]������������������̋�U��EP�MQ�URh��������]����������������̋�U��EPj �MQhw������]������������������̋�U��EP�MQ�URhw������]����������������̋�S�܃������U�k�l$���   �XD3ŉE��C��M��U��U�C��M��U����U��}�w@�E��$� ��E�   �4�E�   �+�E�   �"�E�   ��E�   ��K�   �E�    �}� ��   �U�P�K��Q�U�R��������ul�C�E�}�t�}�t�}�t� �M����M��U������U��C�@�]��	�M�����M��S��R�C��P�KQ�U�R�E�P��p���Q�����h��  �U�P�</����ǅl���    �K�9t�=�Z u�SR�4������l�����l��� u�C�Q��,�����M�3��!����]��[�ȉ�щډȉ��������������������������������������������������������������������������������������������������������������������̋�U����E�]��E�  �E��M���  �U����f�M��E���]��������������������������̋�U��Q�E%�  ��f�E��M����  f�M��E���]��������������������̋�U���E%�  ���ȋU�����P���E�$�Y����]��������������̋�U����E�]��E%�  �M���f�E��E���]����������������������̋�U��}  �u�} u�   �X�}  ��u�} u�   �B�E%�  =�  u�   �+�M���  ���  u�U����u�} t�   �3�]�������������������������������������������̋�U������]����Dz���]��E�    ��   �E%�  ��   �M����u
�} ��   �E�������]����Au	�E�   ��E�    �U�U��E��u/�M��M�U��   �t	�E���E�M��M�U����U����E%��  f�E�}� t�M�� �  f�Mj ���E�$������]��.j ���E�$�t�����]��U���  ����-�  �E��M�U���E���]���������������������������������������������������������������������������������̋�U����E���]��E���]���������̋�U������]��E�E��M������U��   �ʉM��E���]���������������̋�U������]��E�E��M������U�ҁ�   �ʉM��E���]�������������̋�U��EP���E�$�L�����]��������������������̋�U������]�h��  h?  �H*�����E��E%�  =�  ��   ���E�$�~&�����E�}� ~C�}�~�}�t�5h��  �M�Q��)�����E�   �U�R���E�$j%��$�����   �E�P�E�X.���$���E�$j%j��������o���]����Dz)�M�Q��W�����$���E�$j%j�������:�U�R���E�$�d����؃��E����E��E��]�h��  �M�Q�>)�����E���]��������������������������������������������������������������������������������̋�U���0���]�h��  h?  ��(�����E��E%�  =�  t�M���  ���  ��   �U���  ���  u�E����u(�} u"�M���  ���  uC�U����u�} t3�E�P�E�E���$���E�$���E�$j&j�Z�����$�X  �M���  ���  t�U���  ���  u%�E�P���E�$���E�$j&�#�����  �E�]����Dzh��  �M�Q��'�����E��  ���]����Dz$�E�   �E�]����z	�E�    ��E�   ����]����z�E�]����At���]����Au-�E�]����z �U���U��E�E�} u	�M���M��P���]����z�E�]����{���]����Au+�E�]����Au�U���U��E�E�}� u	�M���M��U����  uv�E�����u�}� tf�M�Q���E��$�������]��U��   R���E��$�Z�����]��E�P���E��$���E�$���E�$j&j������$�   �}�  �u�}� t�}�  ��ui�}� uc�M�Q���E��$�6������]ЋU܁�   R���E��$�������]��E�P���E��$���E�$���E�$j&j������$�h��  �M�Q��%�����E���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���E%�  =�  u3���   ]����������������̋�U���E%�  =�  u�M����u�} u�U���  ���  u�   �3�]������������������������������̋�U����E%�  =�  uD���E�$� �����E��}�t�}�t�}�t��   �{�   �t�   �m�   �f�M�� �  �M��U���  u!�E����u�} t�E��������   �,���]����Dz�E���������@��E����%���   ��]����������������������������������������������������������̋�U��Q3��} ���E��}� uh�j j$h��j�^�������u̃}� u-�����    j j$h��hh�h��6�����   ��U�$X�3���]���������������������������������������̋�U��Q3��} ���E��}� uhX�j j-h��j��������u̃}� u-�@���    j j-h��h8�hX�������   ��U�(X�3���]���������������������������������������̋�U��Q3��} ���E��}� uh̊j j6h��j��������u̃}� u-����    j j6h��h��h̊�������   ��U� X�3���]���������������������������������������̋�U����} t�} w�} u�} t	�E�    ��E�   �E��E��}� uh��j j?h��j�Z�������u̃}� u0�����    j j?h��hp�h���2�����   �<  �} t�U� 3��} ���E��}� uh<�j jDh��j���������u̃}� u0�j���    j jDh��hp�h<��������   ��   �} t�}t	�E�    ��E�   �U�U�}� uh��j jEh��j�l�������u̃}� u-�����    j jEh��hp�h���D�����   �Q�M���XR���������M��} u3��,�U�;Ev�"   ��M���XR�EP�MQ�������]��������������������������������������������������������������������������������������������������������������������������������̋�U��$X]����̋�U��(X]����̋�U�� X]����̋�U�츰X]����̋�U��j�h�.h"�d�    P��SVW�XD1E�3�P�E�d�    �=�v uEj�������E�    �=�v u��   ��v����v�E������   �j�&����ËM�d�    Y_^[��]����������������������������������������������̋�U��j�h�.h"�d�    P��SVW�XD1E�3�P�E�d�    j�g������E�    �H   �E������   �j�f%����ËM�d�    Y_^[��]�����������������������������̋�U��j�h�.h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    �E�    �E�    �E�    �E�    �E�    j�������E�    ����E�j h�   h��h��h���E�P������P�������j h�   h��h��hl��M�Q�������P�������j h�   h��h��h4��U�R� ����P����������E���v    �`Y�����`Y�TYh��������Eă}� t�M�����.  �=�v tj��vP��������v    h@v��������   ��v   �@vk�<�M���v��t��vk�<EЉE���v��t$�=�v t�E�   ��v+�vk�<�U���E�    �E�    �E�Pj j?�M܋Rj�hDvj �E�P�ؒ��t�}� u�M܋�B? ��E܋� �U�Rj j?�E܋HQj�h�vj �U�R�ؒ��t�}� u�E܋H�A? �	�U܋B�  �E�   ��   �=�v t#��vQ�U�R�?������u�E�   �   �=�v tj��vP������h  hH�j�M�Q��������P���������v�=�v u	�E�   �Bj h  h��h��h���U�R�E�P�������P��vQ��	����P�\������U�R�������E�P�������M�Q�l�����E������   �j��!����Ã}� ��  j h-  h��h��h��j�U�Rj@�E܋Q�������P��������Uă��UċE����-u�Ũ��ŰEă��EċM�Q�����i�  �EЋU����+t�M����0|�E����9�Uă��U��ԋE����:��   �Uă��UċE�P�)����k�<EЉEЋM����0|�E����9�Uă��U��ߋE����:u<�Uă��UċE�P������EЉEЋM����0|�E����9�Uă��U��߃}� t�E��؉EЋM���Uԃ}� t8j h`  h��h��hP�j�E�Pj@�M܋QR������P�������	�E܋H� �U�R�5������E�P��������M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���	���M�]���������������̋�U���_���M�]���������������̋�U���?����M�]���������������̋�U��j�h�.h"�d�    P���SVW�XD1E�3�P�E�d�    j��������E�    �EP�T   ���E��E������   �j������ËE�M�d�    Y_^[��]��������������������������������̋�U����E�    j h.  h��h�hl��E�P�������P��������}� u3��  �M�Q;TYu�E�H;`Y��  �=�v �G  ��v��uO��vP��vQ��vR��vPj ��vQ��vR��vP�M�QRjj�g  ��,�G��vP��vQ��vR��vP��vQj j ��vR�E�HQj j�  ��,��v��uO��vP��vQ��vR��vPj ��vQ��vR��vP�M�QRjj ��  ��,�G��vP��vQ��vR��vP��vQj j ��vR�E�HQj j �}  ��,�   �E�   �E�   �E�   �E�   �U�zk}�E�   �E�   �E�
   �E�   j j j jj j �E�P�M�Q�U�BPjj�  ��,j j j jj j �M�Q�U�R�E�HQjj ��  ��,�XY;dY}K�E�H;XY|�U�B;dY~3���   �M�Q;XY~�E�H;dY}
�   �   �F�U�B;dY|�M�Q;XY~
�   �   �E�H;dY~�U�B;XY}3��e�M�Qk�<�E�ʋU�Bi�  �i��  �M��M�Q;XYu�E�;\Y|	�   ��3����M�;hY}	�   ��3���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���VW�E�    �}�M  �E%  �yH���@��u�E��d   ����u#�El  ���  ����t�U��Y�E���M���X�U��E����E��M��Fi�m  M��E���������E����d   ��+��E+  ���  ����D1�   ���U�U�;U�E+E�M��k�M�ȉM���U+U�Ek�E�E��}ud�M��  �yI���A��u�E��d   ����u#�El  ���  ����t�U��Y�E���M���X�U�E�;E�~	�M����M��b�U��  �yJ���B��u�E��d   ����u#�El  ���  ����t�U��Y�E���M���X�U�E�E��M�M �M��}u4�U��XY�E$k�<E(k�<E,i��  E0�\Y�M�TY�   �U��dY�E$k�<E(k�<E,i��  E0�hYj h�  h��h@�h4��M�Q������P�������U�i��  hY�hYy �hY \&�hY�dY���dY�+�=hY \&|�hY�� \&�hY�dY���dY�M�`Y_^��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��� V�E�    �E�E�3Ƀ} ���M�}� uhp�j j7hp�j�^�������u̃}� u0������    j j7hp�hT�hp��6������   �u  j$h�   �EP�����3Ƀ} ���M��}� uhDdj j;hp�j���������u̃}� u0�g����    j j;hp�hT�hDd�������   ��  �E��M��P�U�}�� |	�}�@W��s�����    �   ��  �}�| 	�}��&A�v������    �   �  j h�3��E�P�M�Q������F�E�E��F�j h�3�RP�s����M�+ȋE�M��E�E���������E����d   ��+ȋE�+  ���  ���D�j h�Q RP�����M�+ȋE�M��E�}� }|�}� su�M����3��U�� �M��U�E���E�M��  �yI���A��u�E왹d   ����u�E�l  ���  ����u�U��Q �E�� �U��E�M����M��@�U��  �yJ���B��u�E왹d   ����u�E�l  ���  ����u	�U����U��E�M�Hj h�Q �U�R�E�P�$����M�A�U�B�j h�Q RP�����M�+ȋE�M��E�}� t	�E��X��E�Y�E�   �	�M���M�U�E��M��;Q}��E���E�M�U�Q�E�M�U��@+��M�A�Uj h�Q �BP�
Q��������   ���E�Pj h  �M�Q�U�R�\����M�A�U�B�j h  RP�L����M�+ȋE�M��E�j j<�M�Q�U�R� ����M�A�U�Bk�<��M�+ȋE�U�
�E��@     3�^��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����c����E��}� u3�� �EP�M�Q��������E��}� t3���E���]������������������̋�U����E�    �E�E�3Ƀ} ���M�}� uhp�j j7h�j��������u̃}� u0�����    j j7h�h�hp���������   �2  j$h�   �EP�����3Ƀ} ���M�}� uhDdj j:h�j��������u̃}� u0�����    j j:h�h�hDd�n������   �  �E��M�}�@W��}������    �   �  �E��������E��U�iҀ��E�+E�M���F   �U��}�3�|[�E����E��M��3��M�}�3�|=�U����U��E�-�3��E�}� ��|�M����M��U�� ���U��	�E����E��M�U��Q�E����Q ���U�B�E�HiɀQ �U�+щU�}� t	�E��X��E�Y�E�   �	�E����E��M��U��E��;H}��U����U��E�M��H�U�E��M��R+��E�P�M����Q ������   ���E�P�E���  ���U�B�E�Hi�  �U�+щU�E���<   ���U�B�E�Hk�<�U�+ыE��M��A     3���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    ������E��}� u�_����    3��K�E��xD u%h�   h|�jj$�r������M��AD�U��zD t�E��HD�M�������    3���E���]�������������������������������������̋�U��������E��}� u3�� �EP�M�Q�������E��}� t3���E���]������������������̋�U����E�    �E�E�}� |,�}�~�}�t��Di�M��U�Di�y�Di�E��o3�t	�E�   ��E�    �U��U��}� uhX�j j9h��j��������u̃}� u+�����    j j9h��h��hX��W����������E���]���������������������������������������������������̋�U��E�Hi]�����������������̋�U��Hi]����̋�U���<�E�    �e���E��E�    �E�    �E�    �=w ��   hȐ���E؃}� u3���  h���E�P���E�}� u3��  �M�Q�~������wh���U�R��P�a������ whx��E�P��P�D������$wh���M�Q���E�U�R�!������,w�=,w th<��E�P��P��������(w�(w;M�tl�,w;U�ta�(wP�_������Eԋ,wQ�M������EЃ}� t8�}� t2�UԉE�}� t�U�Rj�E�Pj�M�Q�UЅ�t�U���u�E�   �}� t�E    �E�[� w;M�t� wR��������Ẽ}� t�ỦE�}� t,�$w;E�t"�$wQ�������Eȃ}� t
�U�R�UȉE�wP�������Eă}� t�MQ�UR�EP�M�Q�U���3���]������������������������������������������������������������������������������������������������������������������������������������������������̋�U���,�} u�} u�} u3���  �} t�} v	�E�   ��E�    �E�E�}� uh��j jh�j���������u̃}� u0�O����    j jh�hؐh���������   �J  �} u\�U� �}�tI�}���t@�}v:�E��9�Hs��H�M��	�U���U�E�Ph�   �M��Q�/�����3���  �} ��   �U� �}�tI�}���t@�}v:�E��9�Hs��H�M��	�U���U��E�Ph�   �M��Q�������3҃} �U��}� uhЗj jh�j��������u̃}� u0�(����    j jh�hؐhЗ�~������   �#  �M�M��U�U��}�u5�E��M���E���U����U��E���E��t�M����M�t���y�����t&�U;Urh��j j+h�j���������u̋M��U���M���E����E��M���M��t�U����U�t�E���Et�} u�M�� �}� ��   �}�u�UU�B� �P   �?  �E�  �}�tI�}���t@�}v:�M��9�Hs��H�U��	�E���E܋M�Qh�   �U��R�*����������t3�t	�E�   ��E�    �U؉U�}� uhX�j j>h�j���������u̃}� u-�r���� "   j j>h�hؐhX���������"   �p�}�th�}���t_�M+M���;MsQ�U+U����E+�9�Hs��H�M���U+U����E+EԋM�Qh�   �U+U��E�LQ�B�����3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M��1����MQ�UR�EP�MQ�UR�M�����P�*   ���E�M��_����E��]���������������������̋�U��EP�MQ�UR�EP���]�������������������̋�U����EP�M������MQ�UR�EP�MQ�UR�M������P�*   ���E�M�������E��]���������������������̋�U����=4w u3j j jj �����t�4w   ������xu
�4w   �=4wt	�=4w u�EP�MQ�UR�EP����  �=4w�  �E�    �} u�M��B�Ej j �MQ�UR����E��}� u3���   �}� ~63�u2�����3��u���r#h��  �M��T	R�6�����P�F������E���E�    �E��E�}� u3��y�M�Q�U�R�EP�MQ�����u�H�F�} uj j j j j��U�Rj �EP�ؒ�E��!j j �MQ�URj��E�Pj �MQ�ؒ�E��U�R��������E���3���]��������������������������������������������������������������������������������������������������������̋�U��} t�E�M��U���U�E]���������������̋�U��Q�} tV�E���E�M��U��}���  u�EP�%������.�}���  t%3�u!h�j h	  hp�j���������u̋�]��������������������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ���������������������������̋�U��j�h/h"�d�    P���SVW�XD1E�3�P�E�d�    �E������E������}�u!�����     ����� 	   ��������  �} |�E;�ws	�E�   ��E�    �MԉM܃}� uh�fj jNhh�j��������u̃}� u<�=����     �)���� 	   j jNhh�hL�h�f�������������C  �E���M������ x�D
������؉E�uh<fj jOhh�j�)�������u̃}� u<�����     ����� 	   j jOhh�hL�h<f��������������   �UR�.������E�    �E���M������ x�D
��t �MQ�UR�EP�MQ�������E��U��F����� 	   �����     �E������E�����3�uh�ej jZhh�j�N�������u��E������   ��MQ������ËE��U�M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��UR�m������E�}��u;������ 	   3�u!h�ej h�   hh�j�+�������u̃������   �UR�E�P�M�Q�U�R����E��}��u#����E��}� t�E�P�-������������>�M���U������ x�L����U���E������ x�L�E��U���]������������������������������������������������������������������������̋�U��j�h8/h"�d�    P���SVW�XD1E�3�P�E�d�    �}�u�����     �	   �;  �} |�E;�ws	�E�   ��E�    �MԉM��}� uhTj j8h�j��������u̃}� u;�G����     �3���� 	   j j8h�h��hT�������	   �  �E���M������ x�D
������؉E�uhLSj j9h�j�4�������u̃}� u;�����     ����� 	   j j9h�h��hLS�������	   �'  �} |�} r	�E�   ��E�    �UЉU؃}� uh��j j:h�j��������u̃}� u;�6����     �"����    j j:h�h��h���x������   �   �MQ豽�����E�    �U���E������ x�T��t�EP�MQ�UR�������E��43�uh�ej jBh�j���������u������ 	   �E�	   �E������   ��UR�-�����ËE�M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���HV�E�    �E�    �E�    jj j �EP��������E؉U܋M�#M܃��t#jj j �UR��������EЉUԋE�#Eԃ��u�8���� �  �M+MЋUUԉM�U�}� �?  
�}� �3  h   j���P����Eȃ}� u%������    �E�   �E������E�������   h �  �EP�������E�}� |	�}�   r	�E�   ��M�MċUĉU�}� |	�}�   r	�E�   ��E�E��M�Q�U�R�EP��������E�}��u(�T����8u�A����    �E�   �E���E��U��*�E���M�+ȋE�M�E�}� �W���|
�}� �K����M�Q�UR��������E�Pj ���P�`��   �}� ~|�}� svj �MQ�UR�EP�,������E��U��M�#M����tO�UR������P�������؃���E��U��E�#E����u!�n����    �E�   ������]����0�M�#M����t'j �U�R�E�P�MQ�������E��U��U�#U����u	����� �3�^��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�RP�EP��������E��E������]����������̋�U��j�hX/h"�d�    P���SVW�XD1E�3�P�E�d�    �}�u������     ������ 	   ����(  �} |�E;�ws	�E�   ��E�    �MԉM��}� uh�fj jUhȓj��������u̃}� u9�����     �z���� 	   j jUhȓh��h�f�����������  �E���M������ x�D
������؉E�uh<fj jVhȓj�}�������u̃}� u9�����     ������ 	   j jVhȓh��h<f�J���������  ����;U����E�uh��j jWhȓj��������u̃}� u9�����     �����    j jWhȓh��h�������������   �UR�������E�    �E���M������ x�D
��t�MQ�UR�EP��������E��?����� 	   �	����     �E�����3�uh�ej jbhȓj�D�������u��E������   ��EP臶����ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���tV�E������E�E��}�u�ٿ���     ������ 	   ����	  �} |�M;�ws	�E�   ��E�    �U��U��}� u!h�fj h�   hȓj�ܸ������u̃}� u<�g����     �S���� 	   j h�   hȓh��h�f����������y  �M���U������ x�L������ىM�u!h<fj h�   hȓj�P�������u̃}� u<�۾���     ������ 	   j h�   hȓh��h<f�����������  ����;EɃ��M�u!h��j h�   hȓj�۷������u̃}� u<�f����     �R����    j h�   hȓh��h������������x  �E�    �} t �E���M������ x�D
��t3��D  3Ƀ} ���M��}� u!hp�j h�   hȓj�2�������u̃}� u<载���     �����    j h�   hȓh��hp�������������  �E���M������ x�D
$�����E�M�M��}�t�}��  �  �U����҃��U�u!hdUj h�   hȓj聶������u̃}� u<�����     ������    j h�   hȓh��hdU�K���������  �M���s	�E�   ��U��U��E��Eh�   h8�j�MQ�ϯ�����Eԃ}� u�����    胼���    ����  jj j �UR��������M���u������ x�D1(�T1,�   �U����҃��U�u!hdUj h�   hȓj�w�������u̃}� u<�����     ������    j h�   hȓh��hdU�A���������  �M����M�U�UԋEԉEȋM���U������ x�L��H��  �U���E������ x�T��
�r  �} �h  �E���M������ x�EȊL
��Uȃ��UȋẼ��E̋M���M�U���E������ x�D
�U���  �E���M������ x�D
%��
��   �} ��   �M���U������ x�MȊT%��Eȃ��EȋM̃��M̋U���U�E���M������ x�D
%
�E��u{�M���U������ x�L&��
t[�} tU�U���E������ x�UȊD&��Mȃ��MȋŨ��ŰE���E�M���U������ x�D&
j �M�Q�UR�E�P�M���U������ x�Q�ē��t�}� |�U�;Uv^����E܃}�u#����� 	   蝹���M܉�E������  �,�}�mu�E�    �  ��U�R�������E������|  �E�E�E̋M���U������ x�L��   �L  �U����  �}� tE�E����
u:�U���E������ x�T���E���M������ x�T�8�M���U������ x�L����U���E������ x�L�EԉE؋M؉M��U�U�9U��9  �E������   �U���E������ x�T��@u:�E���M������ x�D
���M���U������ x�D��U؋E���
�U؃��U؋E����E��  �  �M����t!�E؋M����E؃��E؋M����M��y  �ŰEԍL�9M�sG�U��B��
u�M����M��U��
�E؃��E���M؋U����M؃��M؋U����U��#  �E����E��E�    j �M�Qj�U�R�E���M������ x�
P�ē��u	����E܃}� u�}� u�M���U؃��U��   �E���M������ x�D
��HtH�M��
u�U��
�E؃��E��,�M���U؃��U؋E���M������ x�E�D
�R�M�;M�u�U��
u�E�� 
�M؃��M��0jj�j��UR��������E��U��E��
t�M���U؃��U������E�+EԉE��M����  �}� ��  �U؃��U؋E����   u�U؃��U��O  �E�   �E����pY��u"�}��E�;E�r�M؃��M؋U����U��͋E����pY�U��}� u����� *   �E������  �E���;E�u�M�M��M���   �U���E������ x�T��H��   �E���M������ x�E؊ �D
�M؃��M؃}�|(�U���E������ x�U؊�T%�E؃��E؃}�u(�M���U������ x�M؊	�L&�U؃��U؋E�+E��E��j�E��ؙRP�MQ�-������E��UċU�+UԉŰE���P�MQ�U�R�E�Pj h��  �ܒ�Ẽ}� u���P�'������E������  �M�+M�3�9M��E���M������ x�T0�M���M��S  �}� tE�U����
u:�M���U������ x�L���U���E������ x�L�8�E���M������ x�D
����M���U������ x�D�UԉU��E��EЋM�M�9M���  �U������   �M���U������ x�L��@u:�U���E������ x�T���E���M������ x�T��M��U�f�f��M����M��UЃ��U��   �  �E����t#�U��E�f�f�
�U����U��EЃ��E���  �M̋UԍD
�9E�sN�M��Q��
u�EЃ��Eй
   �U�f�
�E����E���M��U�f�f��M����M��UЃ��U��  �EЃ��E��E�    j �M�Qj�U�R�E���M������ x�
P�ē��u	����E܃}� u�}� u�   �U�f�
�E����E��  �M���U������ x�L��H��   �U��
u�
   �M�f��U����U��|�E�E��   �U�f�
�E����E��M���U������ x�M��	�L�U����U��E���M������ x�E�� �D
%�M���U������ x�D&
�\�M�;M�u�U��
u�
   �M�f��U����U��5jj�j��EP�������E��U��M��
t�   �E�f��M����M��E����U�+UԉŰE�;Et�M�Q�[������}��u�ỦU���E�E��E�^��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�hx/h"�d�    P���SVW�XD1E�3�P�E�d�    �}�u蝬���     ����� 	   ����  �} |�E;�ws	�E�   ��E�    �M؉M��}� uh�fj jBhДj裥������u̃}� u9�.����     ����� 	   j jBhДh��h�f�p���������/  �E���M������ x�D
������؉E�uh<fj jChДj��������u̃}� u9訫���     ����� 	   j jChДh��h<f����������   �UR�%������E�    �E���M������ x�D
��t�MQ�UR�EP�O������E��?����� 	   �����     �E�����3�uh�ej jNhДj�S�������u��E������   ��EP薠����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP艭�����E��}��u5������ 	   3�uh@�j jlhДj�J�������u̃���   �EPj �MQ�U�R����E��}��u����E���E�    �}� t�E�P�H���������;�M���U������ x�L����U���E������ x�L�E���]���������������������������������������������������������̋�U��j�h�/h"�d�    P���SVW�XD1E�3�P�E�d�    �} @  t-�} �  t$�}   t�}   t�}   t	�E�    ��E�   �EԉE��}� uh�j j7h��j��������u̃}� u.�m����    j j7h��h��h��õ��������  �}�u�9���� 	   ����  �} |�U;�ws	�E�   ��E�    �EЉE܃}� uh�fj j9h��j�S�������u̃}� u.�տ��� 	   j j9h��h��h�f�+���������  �U���E������ x�T������ډU�uh<fj j:h��j�ؠ������u̃}� u.�Z���� 	   j j:h��h��h<f谴��������   �MQ�������E�    �U���E������ x�T��t�EP�MQ��������E��4����� 	   3�uh�ej jEh��j�/�������u��E������E������   ��MQ�k�����ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E���M������ x�D
%�   �E��M���U������ x�L$�����щU��E�E�}�   $�}�   �a  �}� @  tm�}� �  t$�  �}�   �=  �}�   ��   �  �M���U������ x�L������U���E������ x�L�`  �E���M������ x�D
�   �M���U������ x�D�U���E������ x�T$�​E���M������ x�T$��   �M���U������ x�L�ɀ   �U���E������ x�L�E���M������ x�D
$$��M���U������ x�D$�u�U���E������ x�T�ʀ   �E���M������ x�T�M���U������ x�L$�က��U���E������ x�L$�}� u� �  ��}� u	� @  ���   ��]����������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����} @  t�} �  t�}   t	�E�    ��E�   �E��E��}� u!h@�j h�   h��j���������u̃}� u0�v����    j h�   h��h$�h@��ɯ�����   ��URhHw�d�3���]�����������������������������������������������������̋�U��Q3��} ���E��}� u!h��j h�   h��j�;�������u̃}� u0轹���    j h�   h��hܗh���������   ��U�Hw�3���]���������������������������������̋�U��3�]�������̋�U��=�Z u0�EP���E�$�����$���E�$�MQj�5�����$�!������ !   h��  �UR�=������E]���������������������������������̋�U����E�E�]��=�Z u1�EP���E��$���E�$���E�$�MQj訧����$�!�聸��� !   h��  �UR�������E���]����������������������������������̋�S�܃������U�k�l$���   �XD3ŉE��C P�KQ�SR�h�������u)�E�����E��KQ�SR�CP�KQ�S R�E�P�z������KQ�H�������|����=�Z u>��|��� t5�S R���C�$�����$���C�$�CP��|���Q衦����$�%���|���R������h��  �C P�������C�M�3��>�����]��[��������������������������������������������������������������������������̋�S�܃������U�k�l$���   �XD3ŉE��C(P�K Q�SR�(�������u;�E����E��M������M��C�]��S R�CP�KQ�SR�C(P�M�Q�(������SR���������|����=�Z u?��|��� t6�C(P���C �$���C�$���C�$�KQ��|���R�N�����$�%���|���P�j�����h��  �K(Q�R������C �M�3�������]��[�����������������������������������������������������������������������̋�U����E�@    �M�A    �U�B    �E��t�E��  ��M�Q���E�P�M��t�E��  ��U�B���M�A�U��t�E��  ��E�H���U�J�E��t�E��  ��M�Q���E�P�M��t�E��  ��U�B���M�A�U�������������M�Q���ЋE�P�M�����҃������E�H���ʋU�J�E�����Ƀ������U�B�����M�A�U�������������M�Q���ЋE�P�M��� ��҃����E�H���ʋU�J�g����E��E���t�M�Q���E�P�M���t�U�B���M�A�U���t�E�H���U�J�E���t�M�Q���E�P�M��� t�U�B���M�A�U�%   �E�}�   w�}�   t+�}� tI�}�   t.�K�}�   t�@�M����E��1�M�������E���M�������E���M�����E��M���   �U�t5�}�   t�}�   t�1�E����U�
�"�E������U�
��E������U�
�E%�  ���M��� ��ЋE��}  tT�M�Q ���E�P �M�Q ���E�P �M�U��Y�E�H`���U�J`�E�H`���U�J`�E�M��XP�X�U�B ���M�A �U�B �����M�A �U�E� �Z�M�Q`���E�P`�M�Q`�����E�P`�M�U��YP�װ���EPjj �M�Q�|��U�B����t�M�����E��M�Q����t�E�����U�
�E�H����t�U�����M��U�B���t�M����E��M�Q��t�E���ߋU�
�E����M�}�wb�U��$���E���������   �U�
�@�E���������   �U�
�(�E���������   �U�
��E��������U�
�E������M�t�}�t�}�t.�;�U�%����   �M��%�U�%����   �M���U�%�����M��}  t�U�E�@P���M�U�BP���]�}�e�M�5��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�UR������]�����������������������̋�U��j�EP�MQ�UR�EP�MQ�UR�n�����]�����������������������̋�U���D�E���E��M��t �U��tj�������E�����E��  �M��t �U��tj��������E�����E��q  �M���   �U���  j�������E%   �E��}�   w�}�   tW�}� t �}�   tv��   �}�   ��   �   �M�������z��W�]����W���]؋U�E���   �E�������z��W�]��� X���]ЋM�E���Z�U�������z� X�]����W���]ȋE�E���,�M�������z� X�]��� X���]��U�E���E�����E��E  �M���9  �U���-  �E�    �E��t�E�   �M�������D��   �U�R�E��� �$�������]�M��   �M��}�����}�E���.�]��E�   �   ���]�����Au	�E�   ��E�    �U��U��E��f�E��M��f�M��	�U����U��}����}:�E��t�}� u�E�   �M���M�U��t�E�   ��E�M���M�봃}� t�E����]�U�E����E�   �}� t
j�c������E�����E��M��t�U�� tj �@������E����E�3��}� ����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��� �EP�  ���E�}� t^�M�M��U�U�E�E�M�M��U�U�E �E��M$�M�h��  �U(R�ϼ�����E�P��������u�MQ躺�����E��"� h��  �U(R蛼�����EP薺�����E ��]�������������������������������������������������̋�U��Q�E�E��}�t�}�~ �}�~������ !   ��ߩ��� "   ��]��������������������̋�U��Q�E�    �	�E����E��}�}�M��ͨZ;Uu�E��ŬZ���3���]�������������������������������̋�U��Q�E�� t	�E�   �K�M��t	�E�   �:�U��t	�E�   �)�E��t	�E�   ��M��t	�E�   ��E�    �E���]���������������������������������������̋�U��Q��}��E���]��������������̋�U��Q�}����E���]�������������̋�U�����}��E#E�M��U��#��f�E��m��E���]������������������̋�U����E��t
�-�[�]���M��t����-�[�]������U��t
�-�[�]���E��t	�������؛�M�� t���]����]�������������������������̋�U��Q�=Py t�]���E�    �E���]�������������̋�U��j�h�/h"�d�    P���SVW�XD1E�3�P�E�d�    �e�=Py ��   �E��@tp�=�[ tg�E�    �U�E������Q�M���E�}�  �t�}�  �t	�E�    ��E�   �E�Ëe���[    �M�ΈM�U�E�������U�⿉U�U�M�d�    Y_^[��]�������������������������������������������������������̋�U��Q�=Py t�]��e���U���]�����������������̋�U��Q�=Py t�����E��E���?�E���E�    �E���]����������������̋�U��Q�=Py t袱���E��E���?�E��ݒ����E�    �E���]���������������������������̋�U����=Py t8�P����E��E#E�M��#M���E��U������U��U��E�P���������E�    �E���]�������������������������̋�U��Q�����E��E��?E��E��M�Q詅������]����������������������̋�U��jj �EP�MQ��  ��]���������������������̋�U��jj �EPj ��  ��]�������̋�U��jj �EP�MQ�  ��]���������������������̋�U��jj �EPj �|  ��]�������̋�U��jj �EP�MQ�Z  ��]���������������������̋�U��jj �EPj �,  ��]�������̋�U��jh  �EP�MQ�  ��]������������������̋�U��jh  �EPj ��  ��]��������������������̋�U��jh  �EP�MQ�  ��]������������������̋�U��jh  �EPj �y  ��]��������������������̋�U��jh  �EP�MQ�G  ��]������������������̋�U��jh  �EPj �  ��]��������������������̋�U��jhW  �EP�MQ��  ��]������������������̋�U��jhW  �EPj �  ��]��������������������̋�U��jj�EP�MQ�  ��]���������������������̋�U��jj�EPj �\  ��]�������̋�U��jj �EP�MQ�:  ��]���������������������̋�U��jj �EPj �  ��]�������̋�U��jj �EP�MQ��   ��]���������������������̋�U��jj �EPj �   ��]�������̋�U����EP�M��!����M�胂���x t8�M��u����H�y�  u$jj �UR�EP�i   ���E�M��>����E���E�    �M��*����E��]��������������������������������̋�U��j �EP讪����]�����������̋�U��j�h�d�    P���XD3�P�E�d�    �EP�M��R����E�    �M�M�M�要���P�E�L#Mu;�} t�M�舁������   �M�H#U�U���E�    �}� u	�E�    ��E�   �E؉E��E������M��3����E��M�d�    Y��]��������������������������������������������������������������̋�U��Q�} uhpDj j.hؘj�Z�������u̋Pi���Pi�U�U�j:h��jh   ��z�����M��A�U��z t�E��H���U��J�E��@   �%�M��Q���E��P�M����U��J�E��@   �M��U��B��M��A    ��]���������������������������������������������������̋�U����}�u����� 	   3��   �} |�E;�ws	�E�   ��E�    �M��M��}� uh�fj j-hh�j�)�������u̃}� u*諞��� 	   j j-hh�hP�h�f������3��A�=�[�u
�������[�=�[ t�   ��E���M������ x�D
��@��]����������������������������������������������������������������̋�U��j�h0h"�d�    P���SVW�XD1E�3�P�E�d�    3��} ���E؃}� uhmj j6h�j�������u̃}� u.蔝���    j j6h�hܙhm����������   �U�U��޵���� Pj豠�����E�    �ĵ���� P�`������E܋E�Pj �MQ覵���� P�ٵ�����E�蒵���� P�U�R蘘�����E������   ��o����� Pj�]�����ËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������̋�U��Q�E�E��M�Q�UR�EP��v������]������������̋�U��Q�E�E��M�Q�UR�EP辬������]������������̋�U��Q�E�E��M�Qj �UR萬������]��������������̋�U��Q�E�E��M�Q�UR�EP�h�������]������������̋�U��Q�E�E��M�Qj �UR�:�������]��������������̋�U����XD��3�98w���M��} t�XD���U���E�    �E��8w�E���]������������������������̋�U��XD��3�98w����]��������������������̋�U���@�} u�} v�} t	�E�     3���  �} t	�M���������;U����E�uh��j jJh��j��{������u̃}� u0�}����    j jJh��hd�h���ӏ�����   �\  �UR�M�躅���M��{��� �x ��   �M���   ~C�} t�} v�URj �EP�n���������� *   �������M؍M�轚���E���  �} tw3�;U��؉E�uh��j j]h��j�${������u̃}� u=覙��� "   j j]h��hd�h����������E�"   �M��H����E��x  �U�E��} t	�M�   �E�    �M������E��J  �=  �E�    �U�Rj �EP�MQj�URj �M���y��� �HQ�ؒ�E��}� t
�}� ��   �}� ��   �����z��   �} t�} v�URj �EP�&�����3�t	�E�   ��E�    �U��U܃}� uh��j j{h��j��y������u̃}� u:�w���� "   j j{h��hd�h���͍�����E�"   �M������E��L�=���� *   �2�����MȍM�������E��*�} t�U�E���E�    �M��՘���E���M��Ș����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP������]��������������̋�U��� �E������EP�M��Z����M��w��P�MQ�M��w������   P�MQ�U�R豩�����E�}� u�E��E���E������M��M�M��c����E��]�����������������������������������������̋�U����E�����j �EP�Ñ��P�MQ�U�R�/������E��}� u�E��E���E������E��]���������������������̋�U����EP�M��a����M���v����U���   �P�� �  �M�M�薖���E��]����������������������������̋�U��j �EP�|x����]�����������̋�U��EPh  �MQ��}����]�������������������̋�U��h  �EP�ѫ����]�������̋�U��EPj�MQ�}����]������̋�U��j�EP蔫����]����������̋�U��EPj�MQ�S}����]������̋�U��j�EP�T�����]����������̋�U��EPj�MQ�}����]������̋�U��j�EP������]����������̋�U��EPh�   �MQ��|����]�������������������̋�U��h�   �EP�������]�������̋�U��EPj�MQ�|����]������̋�U��j�EP脪����]����������̋�U��EPj�MQ�C|����]������̋�U��j�EP�D�����]����������̋�U��EPh  �MQ� |����]�������������������̋�U��h  �EP������]�������̋�U��EPhW  �MQ�{����]�������������������̋�U��hW  �EP衩����]�������̋�U��EPh  �MQ�`{����]�������������������̋�U��h  �EP�Q�����]�������̋�U��EPj �MQ�{����]������̋�U��j �EP������]����������̋�U���E=�   ���]������������̋�U��Q�EPh  �MQ�z������u�U��_t	�E�    ��E�   �E���]����������������̋�U��Qh  �EP耨������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��Q�EPh  �MQ�z������u�U��_t	�E�    ��E�   �E���]����������������̋�U��Qh  �EP��������u�M��_t	�E�    ��E�   �E���]���������������������S�D$�u�L$�D$3���D$���3��P�ȋ\$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$���؃� [� ������������������������������������������̋�U��=u uj �EP�MQ�URh�W�:   ����j �EP�MQ�URj �   ��]�������������������������̋�U��j�hH�d�    P��H�XD3�P�E�d�    �EP�M��R{���E�    �} t�M�U�3��} ���Ẽ}� uh�j j^h��j�q������u̃}� uD莏���    j j^h��h��h��������E�    �E������M��)����E��  �} t�}|�}$~	�E�    ��E�   �U��Uȃ}� uh0�j j_h��j�vp������u̃}� uD������    j j_h��h��h0��N������E�    �E������M�蓏���E��v  �M�M��E�    �U���E�M����M��M��qo����t0�M��eo������   ~�M��Ro��Pj�E�P�Q������E��j�M�Q�M��.o��P�`i�����E��}� t�U���E�M����M���U��-u�E���E�M���U�E����E���M��+u�U���E�M����M��} |�}t�}$~.�} t�U�E��E�    �E������M�舎���E��k  �>�} u8�M��0t	�E
   �&�U����xt�M����Xu	�E   ��E   �} u8�E��0t	�E
   �&�M����xt�E����Xu	�E   ��E   �}u9�U��0u0�E����xt�U����Xu�M����M��U���E�M����M�����3��u�E�j�U�R�M��m��P��g������t�E��0�E��Qh  �M�Q�M��m��P�g������t0�U��a|�E��z�M�� �M���U�U��E���7�E���f�M�;Mr�\�U���U�E�;E�r�M�;M�u���3��u9U�w�U��UU�U���E���E�} u��M���U�E����E��!����M����M��U��u�} t�E�E��E�    �f�M��u*�U��uV�E��t	�}�   �w�M��u=�}����v4訋��� "   �U��t	�E�������E��t	�E�   ���E�����} t�M�U���E��t�M��ىMЋUЉU��E������M������E��M�d�    Y��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�������]���������������̋�U��=u uj�EP�MQ�URh�W��������j�EP�MQ�URj �n�����]�������������������������̋�U��j�EP�MQ�UR�EP�4�����]���������������̋�U���4  �XD3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M��Pt���E�    3Ƀ} �������������� u!h�nj h  h�Ej�j������u̃����� uF莈���    j h  h�Eh��h�n��}����ǅ��������M��*���������  �E�������������Q��@��   ������P�/������������������t-�������t$������������������� x�������
ǅ����PN�������H$�����х�uV�������t-�������t$������������������� x�������
ǅ����PN�������B$�� ���ȅ�tǅ����    �
ǅ����   ������������������ u!hpmj h  h�Ej�h������u̃����� uF�����    j h  h�Eh��hpm�l|����ǅ��������M�赇��������  3Ƀ} �������������� u!hmj h  h�Ej�h������u̃����� uF葆���    j h  h�Eh��hm��{����ǅ��������M��-���������   ǅ����    �E�    ǅ����    �E�    �E�    �E��������������E���E���  ������ �  �������� |%��������x�������� ����������
ǅ����    ������������������k�	��������@�����������������   3�tǅ����   �
ǅ����    ������������������ u!h�Nj h`  h�Ej�f������u̃����� uF�%����    j h`  h�Eh��h�N�xz����ǅ��������M������������  ��������������������  �������$��1�E�    �M��e��P������R�g��������   ������P�MQ������R�m  ���E��������U���U����������؉�����u!h�Ej h�  h�Ej�e������u̃����� uF�#����    j h�  h�Eh��h�E�vy����ǅ��������M�迄��������  ������R�EP������Q�  ����  �E�    �UԉU؋E؉E�M�M��E�    �E������E�    �  �������������������� ������������wK���������1�$��1�E����E��,�M����M��!�U����U���E��   �E��	�M����M��!  ��������*u(�EP������E�}� }�M����M��U��ډU���E�k�
�������TЉU���  �E�    ��  ��������*u�MQ�~�����EЃ}� }�E�������U�k�
�������LЉM��  ��������������������I������������.�  ���������1�$��1�E���lu�U���U�E�   �E��	�M����M���   �U���6u&�M�Q��4u�E���E�M��� �  �M��   �U���3u#�M�Q��2u�E���E�M�������M��S�U���dt7�M���it,�E���ot!�U���ut�M���xt�E���Xu�ǅ����    ������U��� �U���E�   �E��J
  ��������������������A������������7�  ��������L2�$�2�U���0  u�E�   �E��M���  tUǅ����    �UR�r����f������������Ph   ������Q�U�R�6����������������� t�E�   �&�EP�|����f��|�����|����������E�   �������U��]  �EP�R|������x�����x��� t��x����y u��N�U��E�P�V������E��P�M���   t&��x����B�E���x�����+����E��E�   ��E�    ��x����B�E���x�����U���  �E�%0  u�M���   �M��}��uǅ��������	�UЉ�������������p����MQ�{�����E��U���  te�}� u��N�E��E�   �M���l�����p�����p�������p�����t��l������t��l�������l����ɋ�l���+M����M��[�}� u	��N�U��E���t�����p�����p�������p�����t��t������t��t�������t����ɋ�t���+E��E��  �MQ�z������h�����������   3�tǅ����   �
ǅ����    ��������d�����d��� u!hPEj h�  h�Ej�_������u̃�d��� uF�-~���    j h�  h�Eh��hPE�s����ǅ��������M���~��������  ��  �U��� t��h���f������f����h�����������E�   �  �E�   �������� �������U���@�U��������E��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}У   ~Bh�  hEj�UЁ�]  R�^X�����E��}� t�E��E��MЁ�]  �M���EУ   �U���U�E�H��P���X�����\����M��]��P�E�P�M�Q������R�E�P�M�Q��X���R�TIP��p�����Ѓ��M���   t&�}� u �M��j]��P�U�R�`IP�p�����Ѓ���������gu,�U���   u!�M��3]��P�E�P�\IQ�Zp�����Ѓ��U����-u�M���   �M��U����U��E�P�F������E��	  �M���@�M��E�
   �o�E�
   �f�E�   ǅ����   �
ǅ����'   �E�   �U���   t�E�0��������Q�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�D�������H�����L����   �U���   t�EP��������H�����L����   �M��� tB�U���@t�EP�w��������H�����L�����MQ�w���������H�����L����=�U���@t�EP��v�������H�����L�����MQ��v����3҉�H�����L����E���@t@��L��� 7|	��H��� s,��H����ً�L����� �ډ�@�����D����E�   �E����H�����@�����L�����D����E�% �  u&�M���   u��@�����D����� ��@�����D����}� }	�E�   ��M�����M��}�   ~�E�   ��@����D���u�E�    �E��E��MЋUЃ��UЅ���@����D���t{�E��RP��D���Q��@���R��y����0��T����E��RP��D���P��@���Q�Zw����@�����D�����T���9~��T����������T����E���T�����U����U��g����E�+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@t?�E�%   t�E�-�E�   �(�M���t�E�+�E�   ��U���t�E� �E�   �E�+E�+E䉅<����M���u������R�EP��<���Qj �=	  ��������R�EP�M�Q�U�R�r	  ���E���t$�M���u������R�EP��<���Qj0��  ���}� ��   �}� ��   ǅ$���    �U���8����E܉�4�����4�����4�������4�������   ��8���f�f������������Rj��(���P��0���Q�Ey������$�����8�������8�����$��� u	��0��� uǅ���������&������P�MQ��0���R��(���P�u  ���Z����������Q�UR�E�P�M�Q�S  �������� |$�U���t������P�MQ��<���Rj ��  ���}� tj�E�P��e�����E�    ����������� t������tǅ����    �
ǅ����   �������� ����� ��� u!h�Fj h�  h�Ej�	X������u̃� ��� uC�v���    j h�  h�Eh��h�F��k����ǅ��������M��$w���������������� ����M��w���� ����M�3��{����]Ð�"�#$�$�$�$#%^&a$l$V$K$y$�$ �I �%C&`%N&Y& ��)�&�'�+E'*�&�+�(�+�+�'�+�+�.   	
�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�H��@t�U�z u�E����U�
�p�E�H���U�J�E�x |&�M��E��M���   �M��U����M���UR�EP�e�����E��}��u�M�������U����M���]���������������������������������������������������̋�U��E�M���M��~!�UR�EP�MQ�	������U�:�u���]������������������������̋�U��Q�E�H��@t�U�z u�E�M�U�
�`�E�M���M��~P�U��E��MQ�UR�E�P�������M���M�U�:�u �n���8*u�EP�MQj?�`�������렋�]�����������������������������������̋�U��j�hX0h"�d�    P���SVW�XD1E�3�P�E�d�    �E�����3��} ���E��}� uh�nj j/h؜j�KO������u̃}� u+��m���    j j/h؜hȜh�n�#c��������W�U�B��@t�M�A    �=�UR��������E�    �EP��q�����E��E������   ��MQ�i`����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������̋�U����E�����3��} ���E�}� uhp�j jZh؜j�%N������u̃}� u.�l���    j jZh؜hL�hp���a��������   �U�U��E��H��   ta�U�R�eh�����E��E�P�"Q�����M�Q�O�����P��g������}	�E������$�U��z tj�E��HQ�[�����U��B    �E��@    �E���]�����������������������������������������������������������������������̋�U��j�hx0h"�d�    P���SVW�XD1E�3�P�E�d�    j�'N�����E�    �EP��j����f�E��E������   �j�������f�E�M�d�    Y_^[��]���������������������������������������������̋�U����XD3ŉE�=�[ ts�=�]�u��G���=�]�u���  �   �Pj �E�Pj�MQ��]R����u)�=�[u�����xu��[    ����  �j�
��[   �=�[ uQj j j�E�Pj�MQj �̓P�ؒ�E��=�]�tj �U�R�E�P�M�Q��]R�ȓ��u���  �f�E�M�3���n����]����������������������������������������������������������������������̋�U��j�h�0h"�d�    P���SVW�XD1E�3�P�E�d�    �E�    3��} ���E܃}� u!hp�j h�   h��j��J������u̃}� u<�SQ���     �?i���    j h�   h��h��hp��^��������   �UR��v�����E�j�K�����E�    �E��M����M���t5�Uf�f�EڋM���M�U�R�Dh������=��  u	�E��������E������   �j�k�����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������̋�U���$�} t�} u3���  �E���u�} t3ҋEf�3���  �MQ�M��OS���M��H������   t1�M��H��� ���   th��j jGh �j�
I������u̍M��mH����z u*�} t�Ef��Uf�
�E�   �M��7h���E��R  �M��3H��P�E�Q�3J��������   �M��H������   ~R�M�� H��� �M;��   |=3҃} ��R�EP�M���G������   R�EPj	�M���G����QR�ܒ��uB�M��G��� �M;��   r�U�B��u"�f��� *   �E������M��pg���E��   �M��lG������   �U�M��Mg���E��k�a3��} ��P�MQj�URj	�M��4G��� �HQ�ܒ��u�Af��� *   �E������M���f���E���E�   �M���f���E���M���f����]��������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�b����]�������������������̋�U����EP�M��P���M(Q�U$R�E P�MQ�UR�EP�MQ�UR�M���E��P�.   ��$�E�M���e���E��]�������������������������̋�U���<�=<w u=j j jh��h   j �ԓ��t�<w   ������xu
�<w   �} ~,�EP�MQ��  ���E��U�;U}�E����E��M��M�=<wt�=<w ��  �E�    �E�    �E�    �} u�U��H�M�}$ u�U��H�M$�UR��b�����E��}��u3��  �E�;E$�D  j j �MQ�UR�E�P�M$Q��H�����E��}� u3���  �U��Uj j �EP�MQ�UR�EP�Г�E�}� u�E�    ��   ��   3�u.�}� ~(�}��w"h��  �U��R�q����P�]�����E���E�    �ẺE�}� u�E�    �|�z�M�Qj �U�R�n�����E�P�M�Q�UR�EP�MQ�UR�Г�E�}� u	�E�    �8�E P�MQ�U�R�E�P�M$Q�U�R��G�����E�}� u	�E�    ��E�E�}� t�M�Q�<`�����!�U R�EP�MQ�UR�EP�MQ�Г�E�}� tj�U�R�nQ�����}� t�E;E�tj�M�Q�RQ�����E��e  �=<w�V  �E�    �E�    �E�    �}$ u�U��H�M$j j �UR�EP3Ƀ}( ����   Q�U$R�ܒ�Eԃ}� u3���  �}� ~63�u2�����3��uԃ�r#h��  �MԍT	R��o����P�\�����E���E�    �EȉE؃}� u3��  �M�Q�U�R�EP�MQj�U$R�ܒ��u
�Y  �T  j j �E�P�M�Q�UR�EP�ԓ�E܃}� u
�,  �'  �M��   tI�}  t>�U�;U ~
�	  �  �E P�MQ�U�R�E�P�MQ�UR�ԓ��u
��   ��   ��   �E܉EЃ}� ~63�u2�����3��uЃ�r#h��  �UЍDP��n����P��Z�����E���E�    �MĉM��}� u�|�z�U�R�E�P�M�Q�U�R�EP�MQ�ԓ��u�V�T�}  u+j j j j �U�R�E�Pj �M$Q�ؒ�E܃}� u�'�%�#j j �U R�EP�M�Q�U�Rj �E$P�ؒ�E܃}� t�M�Q�]�����U�R�]�����E���3���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U��E����E���t�M����t�E����E��ۋE+E�����]��������������������������̋�U����EP�M��I���M$Q�U R�EP�MQ�UR�EP�MQ�M���>��P�2   �� �E�M���^���E��]�����������������������������̋�U���$�=@w u8�E�Pjh��j�ܓ��t�@w   ������xu
�@w   �=@wt�=@w ��   �E�    �}  u�M��B�E �} u�M��B�E�M Q�#\�����E�}��u3��  �U�;Ut2j j �EP�MQ�U�R�EP�'B�����E��}� u3��O  �M��M�UR�EP�MQ�UR�E P�ؓ�E��}� tj�M�Q�K�����E��  �=@w�  �E�    �} u�U��H�Mj j �UR�EP3Ƀ}$ ����   Q�UR�ܒ�E�}� u3��   3�u2�}� ~,�}����w#h��  �M�T	R�qj����P�V�����E���E�    �E܉E��}� u3��g�M���Qj �U�R�cg�����E�P�M�Q�UR�EPj�MQ�ܒ�E�}� t�UR�E�P�M�Q�UR�ܓ�E�E�P�EY�����E���3���]�����������������������������������������������������������������������������������������������������������������������������������������������������̋�U���[]����̋�U����&o���E��E��Hl�M��U�;�Wt�E��Hp#�Vu�K���E��U����   ��]�������������������������̋�U��Q�E�x  toj@h�jh�   j�Y�����E��}� u
�   �   �MQ�U�R��   ����t!�E�P�`X����j�M�Q�4I�����   �}�U�ǂ�      ��E� \�E���    \tJ�M���   �´   R�\���u0�E���   ���    h��j jPh@�j�6;������u̋E�M����   3���]����������������������������������������������������������������̋�U����E�    �E�HB�M��U�BD�E��} u�����  �M�M��E�    �U��Rj1�E�Pj�M�Q�%h����E�E�U��Rj2�E�Pj�M�Q�h����E�E�U��Rj3�E�Pj�M�Q��g����E�E�U��Rj4�E�Pj�M�Q��g����E�E�U��Rj5�E�Pj�M�Q�g����E�E�U��Rj6�E�Pj�M�Q�g����E�E�URj7�E�Pj�M�Q�bg����E�E�U�� Rj*�E�Pj�M�Q�Ag����E�E�U��$Rj+�E�Pj�M�Q� g����E�E�U��(Rj,�E�Pj�M�Q��f����E�E�U��,Rj-�E�Pj�M�Q��f����E�E�U��0Rj.�E�Pj�M�Q�f����E�E�U��4Rj/�E�Pj�M�Q�f����E�E�U��Rj0�E�Pj�M�Q�{f����E�E�U��8RjD�E�Pj�M�Q�Zf����E�E�U��<RjE�E�Pj�M�Q�9f����E�E�U��@RjF�E�Pj�M�Q�f����E�E�U��DRjG�E�Pj�M�Q��e����E�E�U��HRjH�E�Pj�M�Q��e����E�E�U��LRjI�E�Pj�M�Q�e����E�E�U��PRjJ�E�Pj�M�Q�e����E�E�U��TRjK�E�Pj�M�Q�se����E�E�U��XRjL�E�Pj�M�Q�Re����E�E�U��\RjM�E�Pj�M�Q�1e����E�E�U��`RjN�E�Pj�M�Q�e����E�E�U��dRjO�E�Pj�M�Q��d����E�E�U��hRj8�E�Pj�M�Q��d����E�E�U��lRj9�E�Pj�M�Q�d����E�E�U��pRj:�E�Pj�M�Q�d����E�E�U��tRj;�E�Pj�M�Q�kd����E�E�U��xRj<�E�Pj�M�Q�Jd����E�E�U��|Rj=�E�Pj�M�Q�)d����E�E�U�   Rj>�E�Pj�M�Q�d����E�E�U�   Rj?�E�Pj�M�Q��c����E�E�U�   Rj@�E�Pj�M�Q�c����E�E�U�   RjA�E�Pj�M�Q�c����E�E�U�   RjB�E�Pj�M�Q�uc����E�E�U�   RjC�E�Pj�M�Q�Qc����E�E�U�   Rj(�E�Pj�M�Q�-c����E�E�U�   Rj)�E�Pj�M�Q�	c����E�E�U�    Rj�E�Pj�M�Q��b����E�E�U�¤   Rj �E�Pj�M�Q��b����E�E�U�¨   Rh  �E�Pj�M�Q�b����E�E�U�°   Rh	  �E�Pj �M�Q�sb����E�E�U�E����   �E��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��} u��  j�E�HQ�@����j�U�BP�@����j�M�QR�y@����j�E�HQ�h@����j�U�BP�W@����j�M�QR�F@����j�E�Q�6@����j�U�B P�%@����j�M�Q$R�@����j�E�H(Q�@����j�U�B,P��?����j�M�Q0R��?����j�E�H4Q��?����j�U�BP�?����j�M�Q8R�?����j�E�H<Q�?����j�U�B@P�?����j�M�QDR�{?����j�E�HHQ�j?����j�U�BLP�Y?����j�M�QPR�H?����j�E�HTQ�7?����j�U�BXP�&?����j�M�Q\R�?����j�E�H`Q�?����j�U�BdP��>����j�M�QhR��>����j�E�HlQ��>����j�U�BpP��>����j�M�QtR�>����j�E�HxQ�>����j�U�B|P�>����j�M���   R�y>����j�E���   Q�e>����j�U���   P�Q>����j�M���   R�=>����j�E���   Q�)>����j�U���   P�>����j�M���   R�>����j�E���   Q��=����j�U���   P��=����j�M���   R��=����j�E���   Q�=����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���VW�E�    �E�    �E�E��E�    �M�y u�U�z ��  jeh�jj0j�AL�����E�}� u
�   �h  �E���   �   �}��jqh�jj�(�����E�}� uj�M�Q�L<�����   �!  �U��    �E�x ��   j}h�jj�Z(�����E��}� u&j�M�Q�<����j�U�R��;�����   ��  �E��     �M�Q>�U��E�Pj�M�Qj�U�R��[����E�E�E��Pj�M�Qj�U�R�[����E�E�E��Pj�M�Qj�U�R�[����E�E�t0�E�P�pC����j�M�Q�[;����j�U�R�M;��������$  �E�HQ��  ���)�E�    �U��\��M��\�Q�E��\�H�U��   �}� t	�E��    ��E�    �E�    �E��\�M���    tA�U���   P�\���u-�M���    w!h��j h�   hH�j�-������u̋E���    t<�M���   R�\���u(j�E���   Q�[:����j�U���   P�G:�����M�U����   �E�M쉈�   �U�E䉂�   3�_^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E���tk�U���0|$�M���9�E���0�U�
�E���E�:�M���;u&�E�E��M��U��B��M����M��U����u��	�M���M닋�]���������������������������������̋�U��} u�[�E�;�\tj�U�P�8�����M�Q;�\tj�E�HQ�s8�����U�B;�\tj�M�QR�T8����]��������������������������������������̋�U���VW�E�    �E�E��E�    �M�y u�U�z �m  jSh�jj0j�G�����E�}� u
�   �  jYh�jj��#�����E��}� uj�E�P�7�����   ��  �M��    �U�z ��  jeh�jj�#�����E�}� u&j�E�P�\7����j�M�Q�N7�����   �  �U��    �E�H8�M��E�    �U��Rj�E�Pj�M�Q�!W����E�E�U��Rj�E�Pj�M�Q� W����E�E�U��Rj�E�Pj�M�Q��V����E�E�U��Rj�E�Pj�M�Q�V����E�E�U��Rj�E�Pj�M�Q�V����E�E�U�� RjP�E�Pj�M�Q�|V����E�E�U��$RjQ�E�Pj�M�Q�[V����E�E�U��(Rj�E�Pj �M�Q�:V����E�E�U��)Rj�E�Pj �M�Q�V����E�E�U��*RjT�E�Pj �M�Q��U����E�E�U��+RjU�E�Pj �M�Q��U����E�E�U��,RjV�E�Pj �M�Q�U����E�E�U��-RjW�E�Pj �M�Q�U����E�E�U��.RjR�E�Pj �M�Q�tU����E�E�U��/RjS�E�Pj �M�Q�SU����E�E�t@�U�R�k=����j�E�P�5����j�M�Q�5����j�U�R�5�����   �>  �E�HQ�a  ����   ��\�}��U���   �M���E���   �U�A�B�M���   �E�J�H�U��   �}� t	�E��    ��E�    �E�    �E��\�M���    tA�U���   P�\���u-�M���    w!h��j h�   hH�j�&������u̋E���    t<�M���   R�\���u(j�E���   Q��3����j�U���   P��3�����M�U䉑�   �E�M����   �U�E艂�   3�_^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E���tk�U���0|$�M���9�E���0�U�
�E���E�:�M���;u&�E�E��M��U��B��M����M��U����u��	�M���M닋�]���������������������������������̋�U��} u��   �E�H;�\tj�U�BP�1�����M�Q;�\tj�E�HQ�1�����U�B;�\tj�M�QR�1�����E�H;�\tj�U�BP�`1�����M�Q; ]tj�E�HQ�A1�����U�B ;]tj�M�Q R�"1�����E�H$;]tj�U�B$P�1����]���������������������������������������������������������������������̋�U���@�XD3ŉE��E�    �E�    �E�    �E�    �E�    �E�E��E�    �M�y ��  �U�z u+�E��Ph  �M�Q0Rj �E�P�TP������t�"  j^h �jj�g�����E�jbh �jjh�  �?�����E�jdh �jjh�  �?�����E�jfh �jjh�  �z?�����E�jhh �jjh  �_?�����E�}� t�}� t�}� t�}� t�}� u�}  �M��    �U�U��E�    �	�E����E��}�   }�M��U���E����E��ۍM�Q�U�BP�����u�&  �}�v�  �M܉Mă}�~S�U�U��	�E����E��M����t8�E��H��t-�U���E��	�M����M��U��B9E��M�M�� ���j j �U�BP�Ḿ�   Qh   �U�Rjj �X���� ��u�  j �E�HQh�   �Uȁ   Rh�   �E��Ph   �M�QRj ��X����$��u�E  j �E�HQh�   �U��   Rh�   �E��Ph   �M�QRj �X����$��u�  3��M�f���   �U��B �E��@ �M�Ɓ�    �U�Ƃ�    �}�~]�E�E��	�M����M��U����tB�M��Q��t7�E���M��	�U����U��E��H9M�� �  �E��M�f��A   ���h�   �Ú�   R�E�P�X)����j�Mȁ�   Q�U�R�@)����j�E�   P�M�Q�))�����U���    ��   �E���   Q�\�����   3�uj j h�   h��j�l������u�j�M���   ���   R��,����j�E���   ��   Q��,����j�U���   -�   P�,����j�M���   R�,�����E��    �M�UЉ��   �E�   �M���   �Ú��   �E���   �Mȁ��   �U���   �E��   �M���   �U�Eĉ��   j�M�Q�,����3���   j�U�R�	,����j�E�P��+����j�M�Q��+����j�U�R��+����j�E�P��+�����   �   �   �M���    tA�U���   P�\���u-�M���    w!hD�j h�   h��j��������u̋Eǀ�       �Mǁ�       ����E���   � ��U���   ����M���   �Uǂ�      3��M�3��	A����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�����N���E��E��Hl�M��U�;�Wt�E��Hp#�Vu�*���E��U����   ��]�������������������������̋�U��Q�} u
�5���E���E����   �U��E���]���������������������̋�U����&N���E��E��Hl�M��U�;�Wt�E��Hp#�Vu�*���E��U��B��]����������������������������̋�U�����M���E��E��Hl�M��U�;�Wt�E��Hp#�Vu�)���E��U��B��]����������������������������̋�U����fM���E��E��Hl�M��U�;�Wt�E��Hp#�Vu�L)���E��E�����]����������������������������̋�U��3�]�������̋�U���(V�E�    �EP�M��)$���M��������   �U��E�    �	�E����E��}�s3�M��U��P�F�������M��U�D�P�F����E��L0�M��jzh��j�U���R�{�����E��}� �  �E��E��E�    �	�M����M��}���   �U��:�E܃��E�j h�   h��hd�h��M��U��P�M����U�+U�+�Q�E�P�Y9����P��#�����M�Q��E����E܉E܋U��:�E܃��E�j h�   h��hd�hx��M��U�D�P�M����U�+U�+�Q�E�P��8����P�#�����M�Q�E����E܉E������U�� �E܃��E܋M��M؍M���7���E�^��]��������������������������������������������������������������������������������������������������������������������������̋�U��j �3����]���������������̋�U���(V�E�    �EP�M���!���M��;������   �U��E�    �	�E����E��}�s4�M��U�D�8P�]D�������M��U�D�hP�HD����E��L0�M��h�   h��j�U���R�'�����E��}� �  �E��E��E�    �	�M����M��}���   �U��:�E܃��E�j h�   h��h$�h���M��U�D�8P�M����U�+U�+�Q�E�P�7����P�!�����M�Q�C����E܉E܋U��:�E܃��E�j h�   h��h$�h8��M��U�D�hP�M����U�+U�+�Q�E�P�6����P�-!�����M�Q�,C����E܉E������U�� �E܃��E܋M��M؍M��5���E�^��]���������������������������������������������������������������������������������������������������������������������̋�U��j � ����]���������������̋�U���,V�E�    �EP�M�����M���������   �U��E�    �	�E����E��}�s3�M��U��P�B�������M��U�D�P��A����E��L0�M���E�    �	�U����U��}�s4�E��M�T�8R��A�������E��M�T�hR�A����E��D0�E�뽋M􋑘   R�A�������E􋈜   Q�{A����E��T0�U��E􋈠   Q�_A�����U��D�E��M􋑤   R�CA�����M��T�U��E􋈨   Q�'A�����U��D�E��M����   �M�h�   h��j�U�R�������E��}� ��  �E��E؋M����   �M�h�   �U�R�E�P�u�����E�    �	�M����M��}���   �U��E؋M܉�j h�   h��h��h���U��E��Q�U�+U��E�+�P�M�Q��3����P�Q�����U�R�P@�����M܍T�U܋E��M؋U܉T�j h�   h��h��h(��E��M�T�R�E�+E��M�+�Q�U�R�]3����P�������E�P��?�����M܍T�U�� ����E�    �	�E����E��}���   �M��U؋E܉D�8j h�   h��h��h���M��U�D�8P�M�+M��U�+�R�E�P��2����P�f�����M�Q�e?�����U܍D�E܋M��U؋E܉D�hj h�   h��h��hP��M��U�D�hP�M�+M��U�+�R�E�P�r2����P������M�Q� ?�����U܍D�E������M؋U܉��   j h�   h��h��h��E􋈘   Q�U�+U��E�+�P�M�Q�
2����P������U�R�>�����M܍T�U܋E؋M܉��   j h�   h��h��h���U􋂜   P�M�+M��U�+�R�E�P�1����P�6�����M�Q�5>�����U܍D�E܋M؋U܉��   j h�   h��h��h ��E􋈠   Q�U�+U��E�+�P�M�Q�D1����P�������U�R��=�����M܍T�U܋E؋M܉��   j h�   h��h��h���U􋂤   P�M�+M��U�+�R�E�P��0����P�p�����M�Q�o=�����U܍D�E܋M؋U܉��   j h�   h��h��hH��E􋈨   Q�U�+U��E�+�P�M�Q�~0����P������U��UԍM��/���E�^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �X5����]���������������̋�U��EPj �MQ�UR�EP�MQ�,
����]�����������̋�U��j j �EP�MQ�UR�EP��	����]�������������̋�U��j �EP�MQ�UR�EP�MQ��	����]�����������̋�U���\�E�    �E�E��MQ�M����3҃} �U؃}� u!hL�j hm  h��j��������u̃}� u@�b,���    j hm  h��h0�hL��!�����E�    �M��-���E���  3Ƀ} ���Mԃ}� u!h�j hn  h��j�g������u̃}� u@��+���    j hn  h��h0�h��<!�����E�    �M��,���E��P  �E�  3Ƀ} ���MЃ}� u!hصj hq  h��j��������u̃}� u@�j+���    j hq  h��h0�hص� �����E�    �M��	,���E���  �} u�M������ ���   �M���U�U��E��E܋M�M��}� ��  �U��E��}� t�}�%t
��   �  3Ƀ} ���M̃}� u!h��j h�  h��j�������u̃}� u@�*���    j h�  h��h0�h���������E�    �M��;+���E��  �E���E�E�    �M���#u�E�   �E���E�M�Q�U�R�E�P�MQ�UR�E�Q�M���
��P��  ����u�}� v�E�   �   �U���U�   �M��
��P�E�Q�������tf�}�v`�U�B��u03�u!h(�j h�  h��j�������u��E�   �Q�%�E�M���E���E�M���M�U����U��E�M���E���E�M���M�U����U��8����}� u*�}� v$�E�  �M+M��M��M���)���E��   �   �U�� �}� u�}� w��(��� "   �q�E�    �}� u!h�j h�  h��j�0
������u̃}� u=�(���    j h�  h��h0�h�������E�    �M��Q)���E���E�    �M��=)���E���M��0)����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���   V�E�E��M����M��}�v��  �U������$�L��M�y |�U�z	�E�   ��E�    �E��E�}� u!h�j h1  h��j�.������u̃}� u0�&���    j h1  h��h�h������3��(  �UR�EP�M�Q�E��Q��  ���  �U�z |�E�x	�E�   ��E�    �M��M��}� u!h�j h:  h��j�������u̃}� u0�	&���    j h:  h��h�h��\����3��  �EP�MQ�U�B�M�T�R�B  ���Y  �E�x |�M�y	�E�   ��E�    �U��U�}� u!hh�j hB  h��j��������u̃}� u0�a%���    j hB  h��h�hh������3���  �MQ�UR�E�H�U�D�8P�  ���  �M�y |�U�z	�E�   ��E�    �E��E�}� u!hh�j hJ  h��j�7������u̃}� u0�$���    j hJ  h��h�hh������3��1  �UR�EP�M�Q�E�L�hQ��  ���	  �}  ��   �UR�EP�MQ�URj�EP��  ����u3���  �M�9 u3���  �U��  �M����E��M����E��MQ�UR�EP�MQj�UR�  ����u3��  �   �EP�MQ�UR�EPj �MQ�]  ����u3��S  �U�: u3��D  �E�� �U����M��U����M��UR�EP�MQ�URj�EP�  ����u3���
  ��
  �M�y|�U�z	�E�   ��E�    �E��E�}� u!hعj h�  h��j�u������u̃}� u0��"���    j h�  h��h�hع�J����3��o
  �U R�EP�MQj�U�BP�  ���H
  �M�y |�U�z	�E�   ��E�    �E��E��}� u!hH�j h�  h��j��������u̃}� u0�P"���    j h�  h��h�hH������3���	  �U R�EP�MQj�U�BP��  ���	  �M�y |�U�z	�E�   ��E�    �E��E܃}� u!hH�j h�  h��j�'������u̃}� u0�!���    j h�  h��h�hH�������3��!	  �U�B��   ���U��}� u�E�   �U R�EP�MQj�U�R�(  ����  �E�x |�M�ym  	�E�   ��E�    �U��U؃}� u!h��j h�  h��j�b������u̃}� u0�� ���    j h�  h��h�h���7����3��\  �M Q�UR�EPj�M�Q��R�{  ���2  �E�x |�M�y	�E�   ��E�    �U��Uԃ}� u!hh�j h�  h��j�������u̃}� u0�: ���    j h�  h��h�hh������3��  �M Q�UR�EPj�M�Q��R��  ���  �E�x |�M�y;	�E�   ��E�    �U��UЃ}� u!h0�j h�  h��j�������u̃}� u0����    j h�  h��h�h0�������3��  �M Q�UR�EPj�M�QR�*  ����  �E�x |�M�y	�E�   ��E�    �U��Ũ}� u!hH�j h�  h��j�g ������u̃}� u0�����    j h�  h��h�hH��<����3��a  �M�y�UR�EP�M���   R�  ����EP�MQ�U���   P�  ���  �M�9 |�U�:;ǅ|���   �
ǅ|���    ��|����Eȃ}� u!h��j h�  h��j��������u̃}� u0����    j h�  h��h�h���l����3��  �U R�EP�MQj�U�P�
  ���k  �M�y |�U�zǅx���   �
ǅx���    ��x����Eă}� u!h�j h�  h��j���������u̃}� u0�j���    j h�  h��h�h������3���  �U�B�E��a  �\  �M�y |�U�zǅt���   �
ǅt���    ��t����E��}� u!h�j h�  h��j�G�������u̃}� u0�����    j h�  h��h�h������3��A  �U R�EP�MQj�U�BP�c	  ���  �M�y |�U�zǅp���   �
ǅp���    ��p����E��}� u!h�j h�  h��j��������u̃}� u0����    j h�  h��h�h��l����3��  �U�z u	�E�   ��E�H���M��U�z |�E�xm  ǅl���   �
ǅl���    ��l����M��}� u!h��j h�  h��j���������u̃}� u0�j���    j h�  h��h�h�������3���  �E�H;M�}	�E�    �-�U�B��   ���E��U�B��   ��;U�|	�U����U��E P�MQ�URj�E�P��  ���}  �}  t+�MQ�UR�EP�MQj�UR�]	  ����u3��S  �)�EP�MQ�UR�EPj �MQ�2	  ����u3��(  �  �UR�EP�MQ�URj�EP�	  ����u3���  ��  �M3҃y �U��}� u!hl�j h  h��j��������u̃}� u0����    j h  h��h�hl��d����3��  �M�A��d   ���U��U R�EP�MQj�U�R�  ���T  �E�x����|�M�y�  ǅh���   �
ǅh���    ��h����U��}� u!hضj h#  h��j���������u̃}� u0�M���    j h#  h��h�hض�����3���   �M�A��d   ���ȃ�k�d�U�B��d   ��ʉM��E P�MQ�URj�E�P��  ���{�����MQ�UR�%���M3҃y  ��P�5  ���O�M��%�E����U�
�E����U�
�+�)3�u!h��j h@  h��j���������u�3���   ^��]ÍI ���>���������'�ԉ%�!��Ď���6�P�`��^�u�O��  	
������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�8 t;�M���t1�E��U���M����E��M���M�U����M��]����������������������̋�U��Q�E�    �} t�EP�MQ�UR�   ���}�E�M;sj�U���U�	�E���E�M��t2�E��
   ����0�E��E��E��
   ���E�U����U�뽋E�M��U�
�E�+M��U�
�	�E�     ��]������������������������������������������������������̋�U����E��M��U�:vE�E��
   ����0�E���M����M��U����M��E��
   ���E�} ~�U�:w��E��M�U�E���M����M��U���E��M��U���M����M��U�E���M���M�U�;U�r̋�]��������������������������������������������������̋�U���X�E�Eȃ}� t�}�t��M���   �U���E���   �M���U���   �E�M���   �?  �}t���U������EЋM�Q��l  f�UԋE�H��f�M֋Uf�Bf�EڋMf�Qf�U܋Ef�Hf�MދUf�f�E�3�f�M�j j �U�R�E�Pj �M���   R�UЉE�}� ��   h��  �E��P�����P�
�����Ẽ}� ��   �M�Q�U�R�E�P�M�Qj �U���   P�UЉE�M̉M��U���U�}� ~9�E�8 v1�M��E���
�U����M��U����U��E����U�
븋E�P�j�����   ��  �M������  �E�8 ��  �E� �E�    �E�    �M�M��	�U����U��E���U���U����U�;�u�܋E����E��M���UċEă�'�Eă}�R�b  �M������$����E��E��M����M��}�w!�U��$�4��E�   �E�m�
�E�b��E�B�  �E��E��M����M��}�w!�U��$�D��E�   �E�d�
�E�a��E�A��  �E��E��}�t�}�t�
�E�y��E�Y�  �M��M��}�t�}�t	��E�   �E�I�  �U��U��}�t�}�t	��E�   �E�H�p  �E��E��}�t�}�t	��E�   �E�M�L  �M��M��}�t�}�t	��E�   �E�S�(  hԼ�U�R�������u�E���E��hм�M�Q�������u	�U���U��E�p��  �E�x�M���   �U���E���   �M��}���   �U�: ��   �EP�M��R�r�������tn�E�8vf�M��Q��u,3�u!h0�j h�  h��j��������u�3��P  �U��M����E����U�
�E����E��M����E��M��E���
�U����M��U����U��E����U�
��   �E������   �U�: ��   �EP�M��R��������tn�E�8vf�M��Q��u,3�u!h0�j h�  h��j���������u�3��}  �U��M����E����U�
�E����E��M����E��M��E���
�U����M��U����U��E����U�
�-����E��E��2����M�����   �U�U��U�E������   �U�: ��   �E����'u�U���U��   �EP�M��R��������tn�E�8vf�M��Q��u,3�u!h��j h�  h��j���������u�3��q  �U��M���E����U�
�E���E�M����E��M��E��
�U����M��U���U�E����U�
�����	�E�E��E��!����M��t;�U�R�EP�MQ�UR�EP�M�Q�UR��������u3���   �E��E��   �MQ�U��P��������tk�M�9vc�U��B��u)3�u!h��j h�  h��j���������u�3��h�E��U���M����E��M���M�U����M��U��M���E����U�
�E���E�M����E��(����   ��]á����a�����B�f�љט�� 







































































	�����������ȘΘ�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����f���E��E��Hl�M��U�;�Wt�E��Hp#�Vu�L����E��]��]������������������������������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^���������������������������̋�U��Q�E�    �} u3��S  �}��   �	�E����E��M��9M���   �U���U�E���E�M�Q���t�E�H��U�B�;�t�M�A��U�J�+���   �U�B���t�M�Q��E�H�;�t�U�B��M�Q�+��   �E�H���t�U�B��M�Q�;�t�E�@��M�Q�+��   �E�H���t�U�B��M�Q�;�t�E�@��M�Q�+��X�����	�E����E��M�;Ms>�U���t�M��E�;�t�U��M�+���E���E�M���M�3���]������������������������������������������������������������������������������������������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�����������������̋�U�������   �E��} u�E�P�\  ���  �M��U��E��@�M��A�U��z t#�E��H���t�E���Pjh ���  ���M��A    �U��: ��   �E�������   �E��x t�M��Q���t�M�Q�O  ����U�R�	  ���E��x uG�M�Qj@h���u  ����t0�U��z t�E��H���t�E�P��  ����M�Q�1	  ���0�U��z t�E��H���t�E�P�  ����M�Q�?  ���U��z u3��N  �} t�E�   �E���E�    �M�Q�U�R�E  ���E��}� t!�}���  t�}���  t�E�P�����u3���   j�M��QR����u3���   �} t&�E�M�f�Qf��E�M�f�Qf�P�Ef�M�f�H�} ��   �U�=  u4j h1  h��hL�h0�h�j@�MQ�����P�N������ j@�URh  �E��HQ�����u3��Bj@�U��@Rh  �E��HQ�����u3��j
j�U�   R�E�P�������   ��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�   �E�    �E�;Eb�}� t\�E�E�+����E��M��U��P�M�R�W �����E�}� u�E��M�T��E���}� }�M����M�	�U����U��3��}� ����]�����������������������������������̋�U��Q�E�Q�����3҃��E�P�M�QR�f����3Ƀ����U�J�E�@    �M�y t	�E�   ��U�P�:  ���E��M�U��Qjh0����E�H��   t�U�B%   t�M�Q��u
�E�@    ��]����������������������������������������������������������̋�U���   �XD3ŉE�����   ��|����EP��  ����x���jx�M�Q��|����B���%���  P��x���Q�����u��|����B    �   �  �E�P��|����QR�n��������r  jx�E�P��|����Q��ҁ������  R��x���P�����u��|����A    �   �G  �U�R��|����Q�	�������u:��|����B  ��|����A��|�����x����B��|�����x����Q��   ��|����H����   ��|����z tt��|����HQ�U�R��|����Q�b�������uQ��|����B����|����A��|�����x����B��|����R��������|���;Au��|�����x����B�E��|����Q��u7��x���P��  ����t$��|����Q����|����P��|�����x����Q��|����H��   ��   ��  jx�U�R��|����H��Ɂ������  Q��x���R�����u��|����@    �   �  �M�Q��|����P�|��������
  ��|����Q��   ��|����P��|����y t7��|����B   ��|����A��|����z u��|�����x����H�   ��|����z tl��|����Q�
������|���;BuP��|���Pj��x���Q�  ����t2��|����B   ��|����A��|����z u��|�����x����H�2��|����B   ��|����A��|����z u��|�����x����H�   ��|����z ut��|����x th�M�Q��|����P�=�������uO��|���Qj ��x���R�c  ����t3��|����H��   ��|����J��|����x u��|�����x����Q��|����@��������M�3��) ����]� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�Q�C����3҃��E�P�M�y t	�E�   ��U�P�!  ���E��M�U��Qjh ����E�H��u
�U�B    ��]��������������������������������������������̋�U���   �XD3ŉE�����   ��|����EP��  ����x���jx�M�Q��|����B���%���  P��x���Q�����u��|����B    �   �  �E�P��|����R��������u`��|����x u��|���Qj��x���R�  ����t3��|�����x����H��|�����x����B��|����Q����|����P�   ��|����y ut��|����z th�E�P��|����R���������uO��|���Pj ��x���Q�  ����t3��|�����x����B��|�����x����Q��|����H����|����J��|����@��������M�3��������]� ������������������������������������������������������������������������������������������������������̋�U��E�HQ�����3҃��E�Pjh�����M�Q��u
�E�@    ]��������������������������̋�U���   �XD3ŉE��9���   ��|����EP�  ����x���jx�M�Q��|����B���%���  P��x���Q�����u��|����B    �   �s�E�P��|����QR�!�������uF��x���P��  ����t3��|�����x����Q��|�����x����H��|����B����|����A��|����B��������M�3�������]� ������������������������������������������������������������������̋�U��E�H��  �U�J���M�A�U�E�H�J]���������������̋�U����XD3ŉE��} t�E���th��UR��������uEj�E�Ph  �M�QR�����u3��ih��E�P�������u����L�M�M�8h ��UR�|������u#j�E�Pj�M�QR�����u3���E�E�MQ��������M�3��������]������������������������������������������������������������������̋�U���f�Ef�E��E�    �	�M����M��}�
s�U��E��E��;�u3���ظ   ��]����������������������̋�U���   �XD3ŉE�V�E%�  �ȁ�   �щ�|���jx�E�Pj��|���Q�����u3��B�U�R�y   ��9Et,�} t&�E�Q�   �����U�P������;�u3���   ^�M�3�������]�������������������������������������������������̋�U����E�    �E��M��U��E���E��tM�M���a|�U���f�E���'�E���M���A|�U���F
�E����E��M����U��DЉE�뚋E���]������������������������������������̋�U����E�    �E��M��U���U�E���A|	�M���Z~�U���a|%�E���z�M����M��U��E��M���M���E���]�������������������������̋�U��Q�} t��}��E�P�V  ���M��} t
��  �U���]��������������������������̋�U�����}��E�P�
  ���E��=Py t�]�M�Q��  ��E���E���]�������������������������������̋�U��QV�}���=Py t�E�P�  �����w  ����M�Q�  ��^��]�������������������������������̋�U����} t^��}��E�P��  ���E�M#M�U��#U�ʉM��E�;E�t'�M�Q�Z  ��f�E��m���}��U�R�  ���E��E�M���} t)�=Py t�UR�EP��  ���M��	�U�    �   ��]��������������������������������������������̋�U��E%����P�MQ�r�����]��������������������̋�U�����}��E�P��  ���E��M#M�U��#U�ʉM�E�;E�t'�M�Q�`  ��f�E��m���}��U�R�  ���E�=Py tB�EP�MQ��  ���E�U�#��E�#�;�t�E�E�   ����E�E����E��]������������������������������������������������̋�U����} 	 u>�}�u8��}��E�%=  ==  u$�=Py t�]��M�����  ���  u�;��7j h[  h��h��h��U������R�EPj ������P���������]��������������������������������������̋�U�������� �E����P����R	  �}� t/�M��Q�%  t �M��Q���U��E��@    �M��A��  ��]�������������������������̋�U����E�    �E��t	�M����M��U��t	�E����E��M��t	�U����U��E��t	�M����M��U�� t	�E����E��M��t�U���   �U��E%   �E��}�   �}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��   �U�t*�}�   t�}�   t�"�E��E���M���   �M���U���   �U��E%   t�M���   �M��E���]��������������������������������������������������������������������������������������̋�U���3�f�E��M��t�U���f�U��E��t�M���f�M��U��t�E���f�E��M��t�U���f�U��E��t�M��� f�M��U��   t�E���f�E��M��   �M��}�   w�}�   t&�}� t�}�   t&�B�}�   t+�7f�U�f�U��-�E�   f�E���M���   f�M���U���   f�U��E%   �E�t�}�   t�}�   t"�(�M���   f�M���U���   f�U��f�E�f�E��M��   t�U���   f�U�f�E���]��������������������������������������������������������������������������������������������������̋�U��Q�E�    �E��?tn�M��t	�U����U��E��t	�M����M��U��t	�E����E��M��t	�U����U��E�� t	�M����M��U��t�E�   �E��E���]�������������������������������������̋�U��Q�����E��E�P�)  ����]������������������̋�U��Q�]��e���U��E�P��  ����]��������������̋�U����E%�E�]��M�Q�   ���E�U#U�E��#E�ЉU��M�;M�u�E��+�U�R��  ���E��E�P��������]��M�Q�2   ����]�������������������������������������������̋�U����E�    �E%�   t	�M����M��U��   t	�E����E��M��   t	�U����U��E%   t	�M����M��U��   t	�E����E��M��   t�U���   �U��E% `  �E��}� @  w�}� @  t$�}� t�}�    t#�:�}� `  t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��@�  �U�}�@t!�}� �  t&�}�@�  t�'�E�   �E���M���   �M���U���   �U��E���]��������������������������������������������������������������������������������������������̋�U����E�    �E��t�M��ɀ   �M��U��t�E�   �E��M��t�U���   �U��E��t�M���   �M��U��t�E�   �E��M��   t�U���   �U��E%   �E��}�   w�}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U��� @  �U���E�    �E���M��� `  �M��U��   �U�}�   t�}�   t�}�   t�$�E�@�  �E���M���@�M���U��� �  �U��E���]��������������������������������������������������������������������������������������������̋�U��Q�E�    �E��?th�M��t	�U����U��E��t	�M����M��U��t	�E����E��M��t	�U����U��E�� t	�M����M��U��t�E�   �E��E���]��������������������������������������������̋�U��Q�E��  �E�P��������]�������������������̋�U��h@]�EP�MQ������]��������������������̋�U���8�E�H
���  ���?  �M�U�B
% �  �E�M�Q�U��E�H�M�U����E�}����u8�E�    �M�Q�I�������t	�E�    ��U�R�������E�   �Z  �E�P�M�Q諼�����U�U܋E�HQ�U�R�n�������t	�E���E�M�U�A+B9E�}�M�Q�Z������E�    �E�   ��   �U�E�;Bk�M�Q�U�R�:������E܉E�M�Q+U�UȋE�P�M�Q�������U�BP�M�Q��������U�B��P�M�Q�������E�    �E�   �~�U�E�;|B�M�Q�������U���   ��U��E�HQ�U�R�O������E��UJ�M��E�   �2�E�M�H�M��U�������U��E�HQ�U�R�������E�    �E�H���    +щU��E��M���E��M���Ɂ�   ���E؋U�z@u�E�M؉H�U�E���M�y u�U�E؉�E���]������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E���E��M����M�E虃�����E�U��  �yJ���B�   +E�   �M���U��E�M��#U�t'�E�P�MQ�_�������u�U�R�EP�L������E�����M���E�M#��E�M���U���U��	�E���E�}�}�M�U��    ��E���]����������������������������������������������������������̋�U����E�������E��E%  �yH���@�   +ȉM����M����҉U��E��M��#U�t3��1�E����E��	�M����M��}�}�U��E�<� t3���߸   ��]��������������������������������������������̋�U����E�������E��E%  �yH���@�   +ȉM�   �M���U�E��M��R�E�P�M��U��P��������E��M����M��	�U����U��}� |)�}� t#�E��M��Rj�E��M��R�������E��ȋE���]������������������������������������������������������̋�U����E�    �EE�E��M�;Mr�U�;Us	�E����E��M�U���E���]����������������̋�U����E�E��M�M��E�    �	�U����U��}�}�E�M����E���E�M����M��Ӌ�]����������������������������������̋�U��Q�E�    �	�E����E��}�}�M��U��    ���]���������������̋�U��Q�E�    �	�E����E��}�}�M��U�<� t3���߸   ��]�����������������������̋�U���V�E�������E��E%  �yH���@�E����M����҉U��E�    �E�    �	�E����E��}�}M�M��U��#E�E�M��U���M���M��U���E��M��U��E��M���    +M�U���U���E�   �	�E����E��}� |.�M�;M�|�U�+U��E��M�u������E��M��    ��^��]������������������������������������������������������������������̋�U��hX]�EP�MQ�������]��������������������̋�U����E�    �E�H
���  f�M��U�B
% �  f�E�M�Q�U�E�H�M��U����E�j@�M�Q��������t�E�   �f�U�f��f�U��E�=�  u�E�   �M�U�Q�E�M���U��E�ЋMf�Q�E���]��������������������������������������������������̋�U���   �XD3ŉEčE��E�3�f�M��E�   �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    3҃}$ �U��}� u!h�j h�   hx�j蓼������u̃}� u0�����    j h�   hx�hP�h��h�����3��  �M�M��U��U��	�E����E��M���� t!�E����	t�U����
t�M����u�Ƀ}�
�s  �E���M��U����U��E���x�����x����G  ��x����$����U���1|�E���9�E�   �M����M��   �U��E$����   ��;�u	�E�   �`�M���t�����t���+t��t���-t#��t���0t�*�E�   �1�E�   3�f�U��"�E�   � �  f�E���E�
   �M����M��  �E�   �U���1|�E���9�E�   �M����M��   �U��E$����   ��;�u	�E�   �j�M���p�����p�����+��p�����p���:w8��p��������$����E�   �+�E�   �"�U����U��E�   ��E�
   �E����E���  �M���1|�U���9�E�   �E����E��K�M��U$����   ��;�u	�E�   �*�E���l�����l���0t�	�E�   ��E�
   �M��M��[  �E�   ��U���E��M����M��U���0|:�E���91�}�s �Mԃ��M��U���0�E���M����M��	�U����U���E��M$����   ��
;�u	�E�   �a�U���h�����h�����+��h�����h���:w/��h�������$� ��E�   �"�E����E��E�   ��E�
   �M����M��w  �E�   �E�   �}� u'��U���E��M����M��U���0u�E����E�����M���U��E����E��M���0|8�U���9/�}�s'�Eԃ��E��M���0�U��
�E����E��M����M���U���d�����d�����+��d�����d���:w/��d�����T��$�H��E�   �"�E����E��E�   ��E�
   �M����M��  �E�   �U���0|�E���9�E�   �M����M���E�
   �U��U��E  �E����E��M���1|�U���9�E�	   �E����E��U�M���`�����`���+t-��`���-t��`���0t�"�E�   �&�E�   �E�������E�   ��E�
   �U��U��  �E�   ��E���M��U����U��E���0u���M���1|�U���9�E�	   �E����E���E�
   �M����M��`  �U���1|�E���9�E�	   �M����M��*�U���\�����\���0t�	�E�   ��E�
   �E��E��  �E�   ǅ|���    ��M���U��E����E��M���0|:�U���91��|���k�
�M��TЉ�|�����|���P  ~ǅ|���Q  �묋�|����E���M���U��E����E��M���0|�U���9���E�
   �E����E��d�}  tN�M����M��U���X�����X���+t��X���-t��E�   �E�������E�   ��E�
   �E��E���E�
   �M����M������U�E���}� �9  �}� �/  �}� �%  �}�v+�M���|	�U����U��E�   �E����E��M����M��}� ��   �U����U��	�E����E��M����u�Eԃ��EԋM����M��ٍU�R�E�P�M�Q�1������}� }�U��ډU��E�E��E��}� u	�M�M�M��}� u	�U�+U�U��}�P  ~	�E�   �B�}�����}	�E�   �0�EP�M�Q�U�R�������f�E�f�E�M��M�U��U�f�E�f�E��3�f�M�3�f�U��E�E؋M؉M�}� u$3�f�U�3�f�E��M�M؋U؉U�E܃��E��V�}� t(��  f�M��E�   ��E�    3�f�U�E܃��E��(�}� t"3�f�M�3�f�U��E�E؋M؉M�U܃��U܋Ef�M�f��U�E�B�M�U؉Q�E��M���Uf�B
�E܋M�3�������]Ë�:����������/����g�t��~�l�u���  �������  �������  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����XD3ŉE���]��`�E��} u�   �} }�M�ىM��^��`�U��} u3��Mf��} tr�U���T�U��E���E�M���M�}� u�׋U�k�U��U�E���� �  |#�U��E�J�M��R�U�E���E�M�M�U�R�EP�������눋M�3��|�����]�����������������������������������������������������������̋�U���L�XD3ŉE�3�f�E��E�    �E�    �E�    �E�    �Mf�Q
f�U�Ef�H
f�M��U��E�3Ё� �  f�U��M���  f�M��UЁ��  f�U��E��M��f�E��U���  }�E�=�  }�M�����  ~2�U���ҁ�   ��� ���E�P�M�A    �U�    �  �E�=�?  "�M�A    �U�B    �E�     ��  �M��u9f�U�f��f�U��E�H�����u�U�z u�E�8 u3ɋUf�J
�  �EЅ�uLf�M�f��f�M��U�B%���u3�M�y u*�U�: u"�E�@    �M�A    �U�    �I  �E�    �E�    �	�E����E��}���   �M���M��E�   �   +U��U��	�Eȃ��Eȃ}� ~x�MM��MċUỦU��E�L؉M��U���M���E��E�P�M�Q�U��P�)������E��}� t�M�f�T�f���E�f�T܋M����M��Ũ��U��y����E���E��<����M����?  f�M��U���~$�E�%   �u�M�Q�w�����f�U�f��f�U����E���Qf�M�f��f�M��U���},�E؃�t	�Mԃ��MԍU�R������f�E�f��f�E��̃}� t�M؃�f�M��U؁� �  �E�%�� = � u_�}��uP�E�    �}��u8�E�    �M����  u� �  f�U�f�E�f��f�E��f�M�f��f�M��	�Uރ��U��	�Eڃ��E��M����  |/�U���ҁ�   ��� ���E�P�M�A    �U�    �-�Ef�M�f��U�E܉B�M�U��Q�E��M���Uf�B
�M�3��K�����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E���   �����ىM��U�B%   �����؉E��M���E��M�Q��U��E�P�M�Q��U��E�P��]������������������������������̋�U����E�H����Ɂ�   ��M��U�B�����%   ��E��M�Q��E�P�M�Q��U��E�P�M���U��E���]���������������������������̋�U����XD3ŉE��EPj j j �MQ�UR�EP�M�Q������ �E�UR�E�P��������E��}�u	�M���M�E�M�3��������]��������������������������������������̋�U���x�XD3ŉE��M  f�E��M   f�M���   f�U��E��C�E���E���E���E���E���E���E���E���E���E���E���E�?�E�   f�Ef�E�M�M؋U�U��E�% �  f�E��M���  f�M��U���t	�E�@-��M�A �U��uM�}� uG�}� uA3��Mf��U��� �  ��҃���-�E�P�M�A�U�B0�E�@ �   �  �M���  �e  �   �Ef��}�   �u�}� tP�M؁�   @uEj j|h��h��hh�h\�j�U��R�������P�~������E�@�E�    ��   �M���tW�}�   �uN�}� uHj h�   h��h��h�h��j�U��R������P�������E�@�E�    �   �}�   �uK�}� uEj h�   h��h��h��h��j�M��Q�9�����P�Ȱ�����U�B�E�    �Cj h�   h��h��hH�h@�j�E��P�������P胰�����M�A�E�    �  �U���f�U��E�%�   f�E��M���f�M��U��E����M��E�����M��E����+U��U��M���f�M�f�U�f�U��E؉E��M��M�3�f�U�j�E���P�M�Q�������U����?  |f�E�f��f�E��M�Q�U�R��������Ef�M�f��U��tP�E�E�E�} @3ɋUf�
�E�- �  �������-�M�A�U�B�E�@0�M�A �   �  �}~�E   �U����?  �U�3�f�E��E�    �	�M���M�}�}�U�R趫������}� },�E���%�   �E��	�M����M��}� ~�U�R�d�������E���E��M���M��	�U���U�}� ~a�E��E̋M��MЋU��UԍE�P�A������M�Q�5������U�R�E�P� ������M�Q�������U���0�E���M����M��E� 됋U����U��E���M�U����U��E��5|[�	�M����M��U��9U�r�E����9u�U��0�ًE��9E�s�M����M��Uf�f���Mf��U���M���k�	�U����U��E��9E�r�M����0u�ߋE��9E�s=3ɋUf�
�E�- �  �������-�M�A�U�B�E�@0�M�A �   �&�U���E�+��M�A�U�B�M�D �E܋M�3�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M�R�E�Q蚪�����E��}� t0�U��Rj�E�HQ�y������E��}� t�U�B���M�A�U��R�E�HQ�U�BP�D������E�}� t�M�Q���E�P�M��Q�U�BP�M�QR��������]�������������������������������������������������̋�U��j
j �EP�)�����]���������̋�U��EPj
j �MQ������]���������������������̋�U��EP�o�����]�������������̋�U��EP�MQ�k�����]���������̋�U��j
j �EP�������]���������̋�U��EPj
j �MQ�M�����]���������������������̋�U����  �XD3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M������E�    3Ƀ} �������������� u!h�nj h  h�Ej�Ϟ������u̃����� uF�N����    j h  h�Ehh�h�n衲����ǅ@��������M�������@����   3��} �������������� u!hmj h  h�Ej�G�������u̃����� uF�Ƽ���    j h  h�Ehh�hm������ǅ<��������M��b�����<����x  ǅ����    �E�    ǅ����    �E�    �E�    �Uf�f�������������U���U���f  ������ �Y  �������� |%��������x�������� �����(����
ǅ(���    ��(���������������k�	��������@�����������������   3�tǅ$���   �
ǅ$���    ��$��������������� u!h�Nj h`  h�Ej�ٜ������u̃����� uF�X����    j h`  h�Ehh�h�N諰����ǅ8��������M��������8����
  �������� ����� ����(  �� ����$����E�   ������Q�UR������P�a  ����  �E�    �MԉM؋U؉U�E�E��E�    �E������E�    ��  ������������������ ����������wL����������$����U����U��-�E����E��"�M����M���U��ʀ   �U��	�E����E��K  ��������*u(�UR�������E�}� }�E����E��M��ىM���U�k�
�������LЉM���  �E�    ��  ��������*u�EP貵�����EЃ}� }�E�������M�k�
�������DЉE��  ������������������I����������.�  ���������$����U���lu�M���M�U���   �U��	�E����E���   �M���6u%�E�H��4u�U���U�E� �  �E��   �M���3u"�E�H��2u�U���U�E�%����E��S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    �w�����M��� �M���U���   �U��t
  ������������������A����������7�P  �������p��$�4��M���0  u	�U��� �U��E�   �EP������f�������M��� tW���������   ������ƅ���� �M�蓘��P�M�芘��� ���   Q������R������P趴������}�E�   �f������f�������������U��E�   �  �EP�S����������������� t�������y u��N�U��E�P�W������E��P�M���   t&�������B�E���������+����E��E�   ��E�    �������B�E���������U���  �E�%0  u	�M��� �M��}��uǅ�������	�UЉ����������������MQ胲�����E��U��� ��   �}� u��N�E��M��������E�    �	�U܃��U܋E�;�����}L���������t?�M�����P�������Q��������t������������������������������d�}� u	��N�M��E�   �U�����������������������������t���������t���������������ɋ�����+U����U��  �EP�}�������|������������   3�tǅ���   �
ǅ���    �������x�����x��� u!hPEj h�  h�Ej苖������u̃�x��� uF�
����    j h�  h�Ehh�hPE�]�����ǅ4��������M�覵����4����  ��  �M��� t��|���f������f����|�����������E�   �  �E�   �������� f�������M���@�M��������U��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}У   ~Ah�  hEj�MЁ�]  Q�:������E��}� t�U��U��E�]  �E���EУ   �M���M�U�B��J���p�����t����M�蓔��P�U�R�E�P������Q�U�R�E�P��p���Q�TIR蟧�����Ѓ��E�%�   t'�}� u!�M��G���P�M�Q�`IR�n������Ѓ���������gu+�M���   u �M�����P�U�R�\IP�7������Ѓ��M����-u�E�   �E��M����M��U�R�$������E��  �E���@�E��E�
   �u�E�
   �l�E�   ǅ����   �
ǅ����'   �E�   �M���   t�0   f�U싅������Qf�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ��������`�����d����   �U���   t�EP���������`�����d����   �M��� tB�U���@t�EP�����������`�����d�����MQ�ڭ���������`�����d����=�U���@t�EP购�������`�����d�����MQ虭����3҉�`�����d����E���@t@��d��� 7|	��`��� s,��`����ً�d����� �ډ�X�����\����E�   �E����`�����X�����d�����\����E�% �  u&�M���   u��X�����\����� ��X�����\����}� }	�E�   ��M�����M��}�   ~�E�   ��X����\���u�E�    �������E��MЋUЃ��UЅ���X����\���t{�E��RP��\���Q��X���R�°����0��l����E��RP��\���P��X���Q�/�����X�����\�����l���9~��l����������l����E���l�����U����U��g���������+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@tN�E�%   t�-   f�M��E�   �2�U���t�+   f�E��E�   ��M���t�    f�U��E�   �E�+E�+E䉅T����M���u������R�EP��T���Qj �P  ��������R�EP�M�Q�U�R�  ���E���t$�M���u������R�EP��T���Qj0�	  ���}� ��   �}� ��   �U���P����E܉�L�����L�����L�������L�����~}�M�莏��P�M�腏��� ���   Q��P���R������P豫������H�����H��� ǅ���������2������Q�UR������P��  ����P����H�����P����j����������R�EP�M�Q�U�R�  �������� |$�E���t������Q�UR��T���Pj �  ���}� tj�M�Q�؜�����E�    �u��������� t������tǅ���    �
ǅ���   �������D�����D��� u!h�Fj h�  h�Ej��������u̃�D��� uC�e����    j h�  h�Ehh�h�F踢����ǅ0��������M�������0������������,����M�������,����M�3�������]Ë�����
��������W�Y�d�N�C�r�{� �I ��;�Y�F�R� ��������D�)������$�����������   	
�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�H��@t�U�z u�E����U�
�4�EP�MQ�|������Ё���  u�E� ������M����E�]����������������������������������̋�U��E�M���M��~!�UR�EP�MQ�Y������U�:�u���]������������������������̋�U��Q�E�H��@t�U�z u�E�M�U�
�b�E�M���M��~R�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u �3����8*u�EP�MQj?��������랋�]�������������������������������������������������̋�U����E�    �E�    �E�H��pt	�U��pu�E�H�U3�;����#  �E�H��st�U�B��St	�E�    ��E�   �M�M��U��st�E��St	�E�    ��E�   �M��M��}� u�}� tA�U�;U�u*�E�H�� ��Ƀ��U�� ��҃�;�u	�E�   ��E�    �E��  �E�H��dtv�U�B��itj�M�Q��ot^�E�H��utR�U�B��xtF�M�Q��Xt:�E��dt1�M��it(�U��ot�E��ut�M��xt�U��X��   �E�H��dtE�U�B��it9�M�Q��ot-�E�H��ut!�U�B��xt�M�Q��Xt	�E�    ��E�   �E��dt6�M��it-�U��ot$�E��ut�M��xt�U��Xt	�E�    ��E�   �E�;E�t3��T�M�Q��   ����ڋE%   �����;�u�M�Q�� ����ڋE�� �����;�t3���M�3�;U����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  �XD3ŉ�X���ǅ<���    ǅ����    ǅ����    ǅp���    ǅ����    ǅx���    ǅ����    �EP��`����؍��ǅ����    ǅ����    ǅH���    ǅ����    ǅ��������ǅ��������ǅ��������ǅ|�������ǅ��������ǅ����    3Ƀ} ����8�����8��� u!h�nj h  h�Ej�:�������u̃�8��� uI蹡���    j h  h�Eh��h�n������ǅ4���������`����R�����4����3  3��} ����4�����4��� u!hmj h  h�Ej诂������u̃�4��� uI�.����    j h  h�Eh��hm聖����ǅ0���������`����ǡ����0����3  ǅT���    �U������ǅH���    ���H�������H�����H�����2  ��H���u������ u�2  ǅ����    ǅ@���    ǅ����    ǅ\���    ǅ��������ǅ����    ǅp���    �������Mǅ��������ǅ��������ǅ|�������ǅ���������Uf�f��L�����L����U���U���C/  ��T��� �6/  ��L����� |%��L�����x��L����� ����������
ǅ����    ��������P�����P���k�	��@�����@�����@�����@�����  �U���%��  �������u\j
������Q�UR藮������~9���������$u+��H��� uh@  j ������R胪����ǅ����   �
ǅ����    �������)  j
������P�MQ�.����������������������U��H��� ��   ������ |#���������$u������d}ǅ����   �
ǅ����    ��������0�����0��� u!h�Nj hP  h�Ej��������u̃�0��� uI�I����    j hP  h�Eh��h�N蜓����ǅ,���������`���������,����,0  ������;�����~��������������������������������������   ��@�����   3�tǅ����   �
ǅ����    ��������,�����,��� u!h�Nj h\  h�Ej��~������u̃�,��� uI�a����    j h\  h�Eh��h�N贒����ǅ(���������`����������(����D/  ��@����������������F,  �������$��9��H��� u	������t��H���u�������u�,  ǅ����   ��T���Q�UR��L���P�=  ����+  ǅt���    ��t�����x�����x���������������������ǅ����    ǅp�������ǅ����    �+  ��L����������������� ������������wj��������:�$��9���������������E���������������4���������������#�������ʀ   ����������������������+  ��L�����*��  ������ u�UR蜗�����������`  j
������P�MQ�ê���������������������U��H��� ��  ������ |#���������$u������d}ǅ����   �
ǅ����    ��������(�����(��� u!h�Mj h�  h�Ej�_|������u̃�(��� uI�ޚ���    j h�  h�Eh��h�M�1�����ǅ$���������`����w�����$�����,  ������;�����~��������������������������������������������������� uG��������Ǆ����   ��������f��L���f���������������������������   ������R��L���Pj��������������R訮��������؉�$���u!h(Mj h�  h�Ej�&{������u̃�$��� uI襙���    j h�  h�Eh��h(M�������ǅ ���������`����>����� ����+  �(  �+���������������� ����� ���P�7����������������� }���������������������ډ������������k�
��L����TЉ������*(  ǅp���    �(  ��L�����*��  ������ u�MQ趔������p����`  j
������R�EP�ݧ��������|������������M��H��� ��  ��|��� |#���������$u������d}ǅ|���   �
ǅ|���    ��|������������� u!hpLj h�  h�Ej�yy������u̃���� uI������    j h�  h�Eh��hpL�K�����ǅ���������`���葘���������)  ��|���;�����~��|�����x������������x�����x�����������|����������� uG��|�����Ǆ����   ��|�����f��L���f��������|������������������   ������Q��L���Rj��|�����������Q�«��������؉����u!h�Kj h�  h�Ej�@x������u̃���� uI迖���    j h�  h�Eh��h�K������ǅ���������`����X���������(  �%  �+��|���������������������R�Q�������p�����p��� }
ǅp����������p���k�
��L����TЉ�p����W%  ��L�����t�����t�����I��t�����t���.�D  ��t�����<:�$�(:�M���lu�E���E��������   �����������������������   �E���6u,�U�B��4u �M���M�������� �  �������   �E���3u)�U�B��2u�M���M������������������d�E���dt7�U���it,�M���ot!�E���ut�U���xt�M���Xu������   �������ǅ@���    ������#�������� ���������������   ��������#  ��L�����p�����p�����A��p�����p���7�H!  ��p������:�$�l:��������0  u�������� ������ǅ����   ������ u�EP�,�����f��D�����  ������ |������d}ǅl���   �
ǅl���    ��l������������� u!hhKj hu  h�Ej�3u������u̃���� uI貓���    j hu  h�Eh��hhK������ǅ���������`����K���������%  ��H��� �  �������������� uG��������Ǆ����   ��������f��L���f���������������������������   ������P��L���Qj��������������P裧��������؉����u!h Jj hy  h�Ej�!t������u̃���� uI蠒���    j hy  h�Eh��h J������ǅ���������`����9���������$  �%  �,������������������������Q�2�����f��D����������� t_��D���%�   �����ƅ��� ��`�����r��P��`�����r������   R�����P��X���Q���������}
ǅx���   �f��D���f��X�����X���������ǅ����   �d  ������ u�MQ胍������ �����  ������ |������d}ǅh���   �
ǅh���    ��h��������������� u!hhKj h�  h�Ej�r������u̃����� uI�
����    j h�  h�Eh��hhK�]�����ǅ���������`���裑���������"  ��H��� �  �������������� uG��������Ǆ����   ��������f��L���f���������������������������   ������Q��L���Rj��������������Q�����������؉�����u!h�Ij h�  h�Ej�yq������u̃����� uI������    j h�  h�Eh��h�I�K�����ǅ���������`���葐���������!  �}  �+��������������������������R芋������ ����� ��� t�� ����x u#��N������������R舝�����������d������%   t/�� ����Q�������� ���� �+���������ǅ����   �(ǅ����    �� ����Q�������� �����������  ��������0  u�������� ��������p����uǅd���������p�����d�����d��������������� u�EP脊������������  ������ |������d}ǅ`���   �
ǅ`���    ��`��������������� u!hhKj h5  h�Ej�o������u̃����� uI�����    j h5  h�Eh��hhK�^�����ǅ���������`���褎���������  ��H��� �  �������������� uG��������Ǆ����   ��������f��L���f���������������������������   ������P��L���Qj��������������P�����������؉�����u!h�Ij h9  h�Ej�zn������u̃����� uI������    j h9  h�Eh��h�I�L�����ǅ ���������`���蒍���� �����  �~  �+��������������������������Q苈������������������ ��   ������ u��N������������������ǅ����    ���������������������;�����}O���������tB��`�����l��P�������Q��n������t������������������������������v������ u��N������ǅ����   ����������������������������������t���������t���������������ɋ�����+��������������-  ������ u�EP�L�������������  ������ |������d}ǅ\���   �
ǅ\���    ��\��������������� u!hhKj h�  h�Ej�Tl������u̃����� uI�ӊ���    j h�  h�Eh��hhK�&�����ǅ����������`����l����������  ��H��� �  �������������� uG��������Ǆ����   ��������f��L���f���������������������������   ������P��L���Qj��������������P�Ğ��������؉�����u!h�Ij h�  h�Ej�Bk������u̃����� uI������    j h�  h�Eh��h�I�����ǅ����������`����Z����������  �F  �+��������������������������Q�S�����������蜡������   3�tǅX���   �
ǅX���    ��X��������������� u!hPEj h�  h�Ej�aj������u̃����� uI������    j h�  h�Eh��hPE�3~����ǅ����������`����y�����������  �e  �������� t������f��T���f����������T����ǅx���   �+  ǅt���   ��L����� f��L�����������@��������������  ��H��� ��  ������ |������d}ǅT���   �
ǅT���    ��T��������������� u!hhKj h�  h�Ej�.i������u̃����� uI譇���    j h�  h�Eh��hhK� }����ǅ����������`����F����������  �������������� uG��������Ǆ����   ��������f��L���f���������������������������   ������R��L���Pj��������������R諛��������؉�����u!h�Hj h�  h�Ej�)h������u̃����� uI訆���    j h�  h�Eh��h�H��{����ǅ����������`����A����������  �-  ��X���������ǅ\���   ��p��� }ǅp���   �7��p��� u��L�����guǅp���   ���p���   ~
ǅp���   ��p����   ~Yh�  hEj��p���]  P�a���������������� t ��������������p�����]  ��\����
ǅp����   ������ u#�E���E�M�Q��A��������������  ������ |������d}ǅP���   �
ǅP���    ��P��������������� u!hhKj h  h�Ej�f������u̃����� uI� ����    j h  h�Eh��hhK�Sz����ǅ����������`���虅����������  ��H���t!h�Hj h  h�Ej�f������u̋����������������������������������������Q��A���������������`����(e��P��t���Q��p���R��L���P��\���Q������R������P�TIQ�(x�����Ѓ���������   t0��p��� u'��`�����d��P������P�`IQ��w�����Ѓ���L�����gu4������%�   u'��`����d��P������Q�\IR�w�����Ѓ����������-u!��������   ��������������������������Q脑�����������  ��������@������ǅ����
   �   ǅ����
   �   ǅp���   ǅ<���   �
ǅ<���'   ǅ����   ������%�   t&�0   f��������<�����Qf������ǅ����   �)ǅ����   ������%�   t��������   �������������� �  �%  ������ u�EP�:�������������������  ������ |������d}ǅL���   �
ǅL���    ��L��������������� u!hhKj h�  h�Ej�kc������u̃����� uI�����    j h�  h�Eh��hhK�=w����ǅ����������`���胂����������  ��H��� �  �������������� uG��������Ǆ����   ��������f��L���f���������������������������   ������P��L���Qj��������������P�ە��������؉�����u!h�Gj h�  h�Ej�Yb������u̃����� uI�؀���    j h�  h�Eh��h�G�+v����ǅ����������`����q����������  �]  �1��������������������������Q�;������������������  ��������   �%  ������ u�EP��������������������  ������ |������d}ǅH���   �
ǅH���    ��H��������������� u!hhKj h�  h�Ej�4a������u̃����� uI����    j h�  h�Eh��hhK�u����ǅ����������`����L����������  ��H��� �  �������������� uG��������Ǆ����   ��������f��L���f���������������������������   ������P��L���Qj��������������P褓��������؉�����u!h@Gj h�  h�Ej�"`������u̃����� uI�~���    j h�  h�Eh��h@G��s����ǅ����������`����:���������  �&  �1��������������������������Q��������������������  �������� �e  ��������@�)  ������ u�MQ��y��������������������  ������ |������d}ǅD���   �
ǅD���    ��D�����|�����|��� u!hhKj h�  h�Ej��^������u̃�|��� uI�n}���    j h�  h�Eh��hhK��r����ǅ����������`����~���������Q  ��H��� �  �������������� uG��������Ǆ����   ��������f��L���f���������������������������   ������Q��L���Rj��������������Q�_���������؉�x���u!h Jj h�  h�Ej��]������u̃�x��� uI�\|���    j h�  h�Eh��h J�q����ǅ����������`�����|���������?  ��  �3����������������t�����t���R��w�������������������(  ������ u!�EP��w���������������������  ������ |������d}ǅ@���   �
ǅ@���    ��@�����p�����p��� u!hhKj h�  h�Ej��\������u̃�p��� uI�C{���    j h�  h�Eh��hhK�p����ǅ����������`�����{���������&  ��H��� �  �������������� uG��������Ǆ����   ��������f��L���f���������������������������   ������P��L���Qj��������������P�4���������؉�l���u!h Jj h�  h�Ej�[������u̃�l��� uI�1z���    j h�  h�Eh��h J�o����ǅ����������`�����z���������  �  �5����������������h�����h���Q��u��������������������Z  ��������@�'  ������ u�EP�u�������������������  ������ |������d}ǅ<���   �
ǅ<���    ��<�����d�����d��� u!hhKj h  h�Ej�Z������u̃�d��� uI�
y���    j h  h�Eh��hhK�]n����ǅ����������`����y����������
  ��H��� �  �������������� uG��������Ǆ����   ��������f��L���f���������������������������   ������P��L���Qj��������������P�����������؉�`���u!h Jj h  h�Ej�yY������u̃�`��� uI��w���    j h  h�Eh��h J�Km����ǅ����������`����x����������	  �}  �2����������������\�����\���Q�s������������������$  ������ u�UR�cs����3ɉ�������������  ������ |������d}ǅ8���   �
ǅ8���    ��8�����X�����X��� u!hhKj h/  h�Ej�cX������u̃�X��� uI��v���    j h/  h�Eh��hhK�5l����ǅ����������`����{w����������  ��H��� �  �������������� uG��������Ǆ����   ��������f��L���f���������������������������   ������Q��L���Rj��������������Q�ӊ��������؉�T���u!h Jj h3  h�Ej�QW������u̃�T��� uI��u���    j h3  h�Eh��h J�#k����ǅ����������`����iv���������  �U  �3����������������P�����P���R�bq����3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�������������������   ��������������������������������������� �  u(������%   u�������������� ��������������p��� }ǅp���   �%�����������������p���   ~
ǅp���   �����������u
ǅ����    ��W�����������p�����p�������p������������������   �������RP������P������Q�St����0�������������RP������R������P�q��������������������9~�������<�������������������������������������K�����W���+���������������������������������   t>������ t���������0t'���������������������0��������������������u��H��� u�]  ��x��� �,  ��������@tj��������   t�-   f������ǅ����   �D��������t�+   f������ǅ����   �!��������t�    f������ǅ����   ������+�����+�������L�����������u��T���Q�UR��L���Pj ��  ����T���Q�UR������P������Q��  ����������t'��������u��T���Q�UR��L���Pj0�y  �������� ��   ������ ��   ��������H�����������D�����D�����D�������D�������   ��`����R��P��`����R������   P��H���Q��D���R�n������@�����@��� ǅT��������2��T���P�MQ��D���R�>  ����H����@�����H����`����!��T���Q�UR������P������Q��  ����T��� |'��������t��T���P�MQ��L���Rj �T  �������� tj������P��_����ǅ����    ������@��� t��@���tǅ4���    �
ǅ4���   ��4�����<�����<��� u!h�Fj h�  h�Ej��Q������u̃�<��� uI�Mp���    j h�  h�Eh��h�F�e����ǅ����������`�����p���������0  �������  ��H��� ��  ǅ����    ���������������������;�������  ����������������0�����0�������0�����0�����   ��0����$��:���������M�������UR�fk�����_  ���������M�������UR�Bk�����;  ���������M�������UR�������  ���������M�������UR�ˀ������   ���������M�������UR��j������   ���������M�������UR�)S�����������������   3�tǅ,���   �
ǅ,���    ��,�����8�����8��� u!h`Fj h-	  h�Ej��O������u̃�8��� uF�An���    j h-	  h�Eh��h`F�c����ǅ����������`�����n���������'�����+�����T�����������`����n����������X���3��r����]ÍI �
�
N����������� �I ���� �D;��$_X^$B�$�$�|$�$o4   	
8B8f8�8�89�8�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�H��@t�U�z u�E����U�
�4�EP�MQ�U�����Ё���  u�E� ������M����E�]����������������������������������̋�U��E�M���M��~!�UR�EP�MQ�Y������U�:�u���]������������������������̋�U��Q�E�H��@t�U�z u�E�M�U�
�b�E�M���M��~R�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u ��]���8*u�EP�MQj?��������랋�]�������������������������������������������������̋�U��j�h�0h"�d�    P���SVW�XD1E�3�P�E�d�    3��} ���E܃}� uhp�j j4h��j�>������u̃}� u-�]���    j j4h��h��hp��jR�������  �M�U�U�E�P�Mt�����E�    �M�Q�UR�S����f�E��E������   ��E�P�O�����f�E��M�d�    Y_^[��]����������������������������������������������������������������������������̋�U���,�XD3ŉE�V�E�H��@�[  �UR�q�������t@�EP�q�������t/�MQ��p���������UR��p��������� x�E���E�PN�E�H$�����у�tj�EP�p�������t@�MQ�p�������t/�UR�p���������EP�p��������� x�E���E�PN�M�Q$������ue�M�Q���E�P�M�y |2�U�f�Mf��U����  f�U�E����U�
f�E��  ��EP�MQ�+d�����  �"  �UR��o�������t@�EP��o�������t/�MQ��o���������UR�o��������� x�E���E�PN�E��H��   ��   �URj�E�P�M�Q��[������t
���  ��   �E�    �	�U����U��E�;E�}m�M�Q���E�P�M�y |.�U��M��T��E�����   �U؋E����U�
��EP�M��T�R��O�����E؃}��u���  �e��E%��  �X�E�H���U�J�E�x |/�M�f�Ef��M����  f�M֋U����M�f�E����UR�EP�b����^�M�3��M^����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EP�MQ��b����]��������̋�U���$h��  h?  �j�����E��E%�  =�  ��   ���E�$��f�����E܃}� ~L�}�~�}�t�>h��  �M�Q�]j�����E�D  �U�R�E���$���E�$j�be�����  �E�P�E�X.���$�E���$���E�$jj�,8����$��  ���]����Dzh��  �M�Q��i�����E��  �U�R���E�$��8�����]�} }!�   �+E9E�}	�E�   ��	�M�M�M������+U9U�~	�E�����	�E�E�E�}� 
  ~G�M�Q���E��$����W�$�d>�����$�E���$���E�$jj�Y7����$�  �}�   ~N�U��   R���E��$��V�����]��E�P���E��$�E���$���E�$jj�7����$�   �}����}6�M�Q�E���.���$�E���$���E�$jj��6����$�   �}����}K�U��   R���E��$�/V�����]��E�P���E��$�E���$���E�$jj�l6����$�,�M�Q���E��$��U�����]�h��  �U�R�h�����E���]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h�0h"�d�    P���SVW�XD1E�3�P�E�d�    3��} ���E��}� uh�j jNh��j�"6������u̃}� u-�T���    j jNh��h��h���I����3��   h�  �UR�G����=�  ��؉E�uh0�j jOh��j�5������u̃}� u*�4T���    j jOh��h��h0��I����3��<j�6�����E�    �UR�k[�����E��E������   �j�m����ËE�M�d�    Y_^[��]������������������������������������������������������������������������������������������������̋�U����8o�E��=y u3���   �}� u"�=@o t�]-����t3���   �8o�M��}� ��   �} ��   �UR�/a�����E��E��8 ��   �M��R�a����;E�v{�E���U����=uj�M�Q�UR�E��Q�	C������uPh�  �U���M��TR��E����=�  r!h@�j h�   h��j��3������u̋M���E��D��M����M��X���3���]�����������������������������������������������������������������������̋�U��j�h�0h"�d�    P���SVW�XD1E�3�P�E�d�    j�w4�����E�    �EP�MQ�UR�EP�X   ���E��E������   �j�`k����ËE�M�d�    Y_^[��]������������������������������������̋�U���3��} ���E��}� u!h��j h�   h��j�2������u̃}� u3�Q���    j h�   h��h��h���^F�����   �   �U�    �} t�} w�} u�} t	�E�    ��E�   �E��E�}� u!h�j h�   h��j��1������u̃}� u3�tP���    j h�   h��h��h���E�����   �   �} t�U� �EP�W�����E��}� u3��d�M�Q�K^�������U��} u3��F�E�;Mv�"   �5j h�   h��h��h���U�R�EP�MQ�[Q����P��;����3���]��������������������������������������������������������������������������������������������������������̋�U��j j j�EP�MQ�UR�G����]���������������̋�U��j�h1h"�d�    P���SVW�XD1E�3�P�E�d�    j�1�����E�    �EP�MQ�UR�EP�MQ�UR�`   ���E��E������   �j�xh����ËE�M�d�    Y_^[��]��������������������������������������������̋�U���3��} ���E�}� u!h��j hX  h��j�/������u̃}� u3�N���    j hX  h��h��h���nC�����   �2  �U�    �} t	�E�     3Ƀ} ���M��}� u!hx�j h^  h��j�/������u̃}� u3�M���    j h^  h��h��hx���B�����   �   �EP��T�����E��}� u3��   �M�Q�w[�������E��UR�EP�MQj�U�R��K�����M��U�: u�M���    �M��� �Ej hr  h��h��h0��E�P�M�Q�U�P�gN����P��8�����} t�M�U��3���]����������������������������������������������������������������������������������������������������������������������̋�U��j�h81h"�d�    P���SVW�XD1E�3�P�E�d�    �d���� �E�3��} ���E؃}� uhmj j4h�j�G-������u̃}� u+��K���    j j4h�h��hm�A��������i�U�R�
c�����E�    �E�P�U�����E܋MQ�UR�EP�M�Q�U���E��U�R�E�P��F�����E������   ��M�Q�S>����ËE��M�d�    Y_^[��]�����������������������������������������������������������������������̋�U��EP�MQ�URh[��"S����]����������������̋�U��EP�MQ�URh����R����]����������������̋�U��EP�MQ�URh����R����]����������������̋�U��EPj �MQh[��R����]������������������̋�U��EPj �MQh���dR����]������������������̋�U��EPj �MQh���4R����]������������������̋�U����E=��  u3�f�M��}�U��   }�E��[�A�E#�f�U��W�MQ�M���4���M��J*����BP�M��<*����QR�E�Pj�MQj�M��"*��P�b������u3�f�U��M���I���E��M#���]������������������������������������������̋�U��Q�E=��  u3��n�M��   }�U��[�P�M#��M�=u u0��VR��VP�M�Qj�URjh�W��a������u3�f�E�j �MQ�UR��0������]�����������������������������������������̋�U���EP�MQ��^����]�������̋�U��} uh�j j0h��j�k)������u̋M�Q��   tK�E�H��t@j�U�BP��6�����M�Q�������E�P�M�    �U�B    �E�@    ]��������������������������������������������̋�U��j j jj jh   �h,��@��|]]����������̋�U��j j jj jh   @h4��@���]]����������̋�U��=�]�t�=�]�t��]P����=|]�t�=|]�t�|]Q���]����������������������������̋�U����XD3ŉE��E� j�E�Ph  �MQ�����u	�E�������U�R�lE�����E��E��M�3��IK����]������������������������̋�U���0�XD3ŉE��E�    �E��M��E�    �U;U��  �E�    �E�P�MQ�����t%�}�u�U�R�EP�����t�}�u�E�   �}� t �}��t�M��M���UR��S�������E��}� u(j j �E�P�MQj�UR�ܒ�E��}� u3��n  3�u2�}� ~,�}����w#h��  �M��T	R�S����P�?�����E���E�    �EЉE�}� u3��  �M���Qj �U�R�}P�����E�P�M�Q�U�R�EPj�MQ�ܒ����   �} t/j j �UR�EP�M�Q�U�Rj �EP�ؒ��t�M�M��   �}� u%j j j j �U�R�E�Pj �MQ�ؒ�E��}� tqh�   h@�j�U�Rj�C�����E��}� tNj j �E�P�M�Q�U�R�E�Pj �MQ�ؒ�E��}� uj�U�R�43�����E�    ��}��t�E�M���}� t�U�R�A�����E��M�3���H����]��������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���8�EP�M���.��3Ƀ} ���M�}� uh�cj j4h��j�$������u̃}� u=�C���    j j4h��h|�h�c�h8�����E�����M��C���E��  3��} ���E��}� uh�bj j5h��j�$������u̃}� u=�B���    j j5h��h|�h�b��7�����E�����M��AC���E��   �M��=#����z u"�EP�MQ��N�����EԍM��C���E��x�b�U��E̍M��#��P�M�Q�?O�����E��U���U�E��MȍM���"��P�U�R�O�����E��E���E�}� t�M�;M�t��U�+U��UЍM��B���EЋ�]����������������������������������������������������������������������������������������������������������̋�U����E��M��U��E���E��A|�}�Z	�M��� �M��U��E��M��U���U��A|�}�Z	�E��� �E��}� t�M�;M�t��E�+E���]������������������������������̋�U����=u ��   3��} ���E��}� uh�cj jbh��j��!������u̃}� u0�q@���    j jbh��h�h�c��5���������   3҃} �U��}� uh�bj jch��j�!������u̃}� u-�@���    j jch��h�h�b�a5���������&�MQ�UR�~L������j �EP�MQ�X������]������������������������������������������������������������������������̋�U���@�} �!  �EP�M���*��3Ƀ} ���M�}� uh�cj j;hp�j� ������u̃}� u=�?���    j j;hp�hP�h�c�n4�����E�����M��?���E��  3��} ���E��}� uh�bj j<hp�j�# ������u̃}� u=�>���    j j<hp�hP�h�b��3�����E�����M��G?���E��1  ����;U����E�uh(�j j=hp�j�������u̃}� u=�2>���    j j=hp�hP�h(��3�����E�����M���>���E��   �M�������z u)�EP�MQ�UR�{�����E̍M��>���E��   �m�E��MčM����P�U�R��J�����E��E���E�M��U��M��d��P�E�P�J�����E��M���M�U���Ut�}� t�E�;E�t��M�+M��MȍM��>���E��3���]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����=u �Y  3��} ���E��}� u!h�cj h�   hp�j��������u̃}� u3�N<���    j h�   hp�h��h�c�1���������  3҃} �U��}� u!h�bj h�   hp�j�`������u̃}� u3��;���    j h�   hp�h��h�b�51���������   ����;M҃��U�u!h(�j h�   hp�j��������u̃}� u0�v;���    j h�   hp�h��h(���0���������.�MQ�UR�EP��������j �MQ�UR�EP�[������]��������������������������������������������������������������������������������������������������������̋�U����XD3ŉE��N@  f�E��M�    �U�B    �E�@    ��M���M�U���U�} vt�E��M�P�U��@�E�MQ�#�����UR��"�����E�P�MQ�������UR��"�����E��M��E�    �E�    �U�R�EP������t����M�y uB�U�B���M�A�U�B���M���M�A�U����M��U���f�U�뵋E�H�� �  u�UR�K"����f�E�f��f�E��؋Mf�U�f�Q
�M�3��O>����]����������������������������������������������������������������������������������������������̋�U��=u uj �EP�MQ�URh�W�:   ����j �EP�MQ�URj �   ��]�������������������������̋�U��j�hx�d�    P��lVW�XD3�P�E�d�    �EP�M���#���E�    �} t�M�U�3��} ���E��}� uh�j j^h�j�������u̃}� uN�8���    j j^h�h �h��r-�����E�    �E�    �E������M��8���E��U��<  �} t�}|�}$~	�E�    ��E�   �U��U��}� uh0�j j_h�j��������u̃}� uN�|7���    j j_h�h �h0���,�����E�    �E�    �E������M��8���E��U��  �M�M��E�    �E�    �U���E�M����M��M�������t0�M���������   ~�M�����Pj�E�P��.�����E��j�M�Q�M����P�������E��}� t�U���E�M����M���U��-u�E���E�M���U�E����E���M��+u�U���E�M����M��} u8�U��0t	�E
   �&�E����xt�U����Xu	�E   ��E   �}u9�M��0u0�U����xt�M����Xu�E����E��M���U�E����E��E�RPj�j��3���E�U�j�M�Q�M����P��������t�U��0�U��Th  �E�P�M��q��P�������t0�M��a|�U��z�E�� �E���M�M��U���7�U���   �E�;Er�   �M���M�U�;U�rLw�E�;E�rB�M�;M�u^�U�;U�uV�u�3��E�RPj�j��K5���u��}��E��U��E�;E�w.r�M�;M�w$�E�RP�U�R�E�P����M�3��։EĉU���U���U�} u��E���M�U����U�������E����E��M��u�} t�U�U��E�    �E�    �   �E��u:�M��u{�U��t�}�   �w!r�}� w�E��uZ�}����rQw�}��vI�%4��� "   �M��t�E������E������&�U��t�E�    �E�   ���E������E�����} t�E�M���U��t�E��؋Mȃ� �ىEĉMȋUĉU��EȉE��E������M��o4���E��U��M�d�    Y_^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�t�����]���������������̋�U��=u uj�EP�MQ�URh�W�:�������j�EP�MQ�URj ������]�������������������������̋�U��j�EP�MQ�UR�EP�������]���������������̋�U��=u uj �EP�MQ�URh�W�:   ����j �EP�MQ�URj �   ��]�������������������������̋�U��j�h��d�    P��@�XD3�P�E�d�    �EP�M��R���E�    �} t�M�U�3��} ���Ẽ}� uh�j jah��j�������u̃}� uD�0���    j jah��h��h���%�����E�    �E������M��)1���E��^  �} t�}|�}$~	�E�    ��E�   �U��Uȃ}� uh0�j jbh��j�v������u̃}� uD��/���    j jbh��h��h0��N%�����E�    �E������M��0���E���  �M�M��E�    �U�f�f�E�M����M��M��o��Pj�U�R��������t�E�f�f�M�U����U����E��-u�M���M�U�f�f�E�M����M���U��+u�E�f�f�M�U����U��} u@�E�P�8������t	�E
   �&�M����xt�E����Xu	�E   ��E   �}uC�U�R��7������u2�E����xt�U����Xu�M����M��U�f�f�E�M����M�����3��u�E��U�R�{7�����E�}��t�V�E��A|	�M��Z~�U��a|9�E��z0�M��a|�U��z�E�� �E���M�M��U���7�U���h�E�;Er�^�M���M�U�;U�r�E�;E�u���3��u9U�w�M��MM�M���U���U�} u��E�f�f�M�U����U��*����E����E��M��u�} t�U�U��E�    �f�E��u*�M��uV�U��t	�}�   �w�E��u=�}����v4�V-��� "   �M��t	�E�������U��t	�E�   ���E�����} t�E�M���U��t�E��؉EЋMЉM��E������M���-���E��M�d�    Y��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP������]���������������̋�U��=u uj�EP�MQ�URh�W�j�������j�EP�MQ�URj �N�����]�������������������������̋�U��j�EP�MQ�UR�EP������]���������������̋�U��� �} uhpDj jdh�Cj�X������u̋M�M��U�R��?�����E��E��H��   u&�*��� 	   �U��B�� �M��A���  �c  �/�U��B��@t$�*��� "   �M��Q�� �E��P���  �2  �M��Q��tJ�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J���  ��  �E��H���U��J�E��H���U��J�E��@    �E�    �M��M�U��B%  u6�OB���� 9E�t�BB����@9E�u�M�Q� ������u�U�R�C�����E��H��  �  �U��E��
+Hy!h`Cj h�   h�Cj��
������u̋E��M��+Q�U��E��H���U��
�E��H���U��J�}� ~�E�P�M��QR�E�P�H3�����E��s�}��t!�}��t�M����U������ x�U���E�PN�E��H�� t9jj j �U�R�I;�����E��U�E�#E���u�M��Q�� �E��P���  �e�M����  �U��Bf��+�E�   �M����  f�M�U�R�E�P�M�Q�2�����E�U�;U�t�E��H�� �U��J���  ��E%��  ��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�    ��E����E��M���M�U�;Us�E���t�ڋE���]��������������������̋�U���<�EP�M�����} u�E�    �M���'���E��  3Ƀ} ���M�}� uh��j j=hx�j�C������u̃}� u=��&���    j j=hx�hP�h��������E�����M��g'���E��  3��} ���E�}� uh4�j j>hx�j��������u̃}� u=�R&���    j j>hx�hP�h4�������E�����M���&���E��!  ����;U����E�uh�j j?hx�j�]������u̃}� u=��%���    j j?hx�hP�h��5�����E�����M��&���E��   �M��}���P�z u(�EP�MQ�UR�EP�f�����E̍M��E&���E��u�M��D���H�QR�EP�MQ�UR�EPh  �M�� ���H�QR�M����P�1���� �E��}� u�E�����M���%���E���E����EčM���%���Eċ�]����������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�l����]�������������������̋�U����E�    �@o�E��M��9 ��   j j j j j��U��Pj j �ؒ�E�}� u����   j=h�jj�M�Q�l"�����E��}� u����rj j �U�R�E�Pj��M��Rj j �ؒ��uj�E�P���������=j �M�Q�F$������}�}� tj�U�R�^�����E�    �E����E��4���3���]�����������������������������������������������������������������������̋�U����EP�M��a���M Q�UR�EP�MQ�UR�EP�M����P�6   ���E�M��#���E��]���������������������������������̋�U��}�}3���EP�MQ�UR�EP�ܓ]����������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��������������������������������̋�U���E��0}����
  �M��:}�E��0��  �U���  ��  �E=`  }�����  �M��j  }�E-`  �  �U���  }����  �E=�  }�E-�  �  �M��f	  }����w  �U��p	  }�E-f	  �]  �E=�	  }����J  �M���	  }�E-�	  �0  �U��f
  }����  �E=p
  }�E-f
  �  �M���
  }�����  �U���
  }�E-�
  ��  �E=f  }�����  �M��p  }�E-f  �  �U��f  }����  �E=p  }�E-f  �{  �M���  }����g  �U���  }�E-�  �M  �E=f  }����:  �M��p  }�E-f  �   �U��P  }����  �E=Z  }�E-P  ��   �M���  }�����   �U���  }�E-�  ��   �E=   }����   �M��*  }�E-   �   �U��@  }����   �E=J  }�E-@  �n�M���  }����]�U���  }�E-�  �F�E=  }����6�M��  }�E-  ������U���  }�E-�  ����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M��Q	���M$Q�U R�EP�MQ�UR�EP�MQ�M�����P�2   �� �E�M��w���E��]�����������������������������̋�U���H�XD3ŉEԃ=Lw u=jh��jh��j j �����t�Lw   ������xu
�Lw   �} ~�EP�MQ��  ���E��}�}3��v  �}  ~�U R�EP�  ���E ��} �}3��N  �=Lwt�=Lw �  �E�    �E�    �} u�M��B�E�}$ u�M��B�E$�MQ�m�����E��}��u3���  �U�;U$trj j �EP�MQ�U�R�E$P�q�����E��}� u3��  j j �M Q�UR�E�P�M$Q�E�����E��}� uj�U�R�����3��~  �E��E�M��M�U R�EP�MQ�UR�EP�MQ����E�}� tj�U�R��
����j�E�P�
�����E��'  �=Lw�  �E�    �}$ u�M��B�E$�} t
�}  �j  �M;M u
�   ��  �} ~
�   ��  �}~
�   ��  �U�R�E$P�����u3��  �} u�} t-�}u�}  t!h��j h�   hH�j�l�������u̃} ~m�}�s
�   �X  �UƉU��	�E؃��E؋M����t8�E��H��t-�U��M��;�|�E��U��B;�
�   �  뵸   ��  �}  ~m�}�s
�   ��  �MƉM��	�U؃��U؋E����t8�U��B��t-�M��E��;�|�U��M��Q;�
�   �  뵸   �  j j �EP�MQj	�U$R�ܒ�E�}� u3��`  �}� ~63�u2�����3��u��r#h��  �M�T	R��'����P������E���E�    �E��E��}� u3��
  �M�Q�U�R�EP�MQj�U$R�ܒ��u
��   ��   j j �E P�MQj	�U$R�ܒ�E܃}� u
�   �   �}� ~63�u2�����3��u܃�r#h��  �M܍T	R�M'����P�]�����E���E�    �E��E�}� u�O�M�M�Q�U�R�E P�MQj�U$R�ܒ��t!�E�P�M�Q�U�R�E�P�MQ�UR����E�E�P�2�����M�Q�&�����E���3��M�3��m����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U��E����E���t�M����t�E����E��ۋE+E�����]��������������������������̋�U���<�EP�M��1���} u�E�    �M��z���E��  3Ƀ} ���M�}� uh�j j?h��j���������u̃}� u=�e���    j j?h��ht�h�������E�����M�����E��  3��} ���E�}� uhL�j j@h��j�p�������u̃}� u=�����    j j@h��ht�hL��H�����E�����M�����E��.  ����;U����E�uh(�j jAh��j���������u̃}� u=����    j jAh��ht�h(���
�����E�����M��!���E��   �M�������z u-�M�����P�EP�MQ�UR�X������E̍M������E��~�M������� �HQ�UR�EP�MQ�URh  �M������ �HQ�M�����P�F!���� �E��}� u����    �E�����M��w���E���U����UčM��a���Eċ�]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��=u u�EP�MQ�UR�3������j �EP�MQ�UR������]������������������̋�U���$V�E�    �E�    3��} ���E܃}� uhl�j jYh��j���������u̃}� u.�O���    j jYh��h��hl����������T  �U��E�}� tj=�M�Q�K%�����E��}� t�U�;U�u�����    ����  �E�+E�=�  |h��j jkh��j�.�������u�h�  �U���R������=�  rh8�j jlh��j���������u̋M��Q��҃��U�8o;<ou�8oQ�g  ���8o�=8o ��   �} t*�=@o t!�_�����t�&���    ����F  �   �}� t3��4  �   �=8o u8h�   h��jj�������8o�=8o u�����  �8o�    �=@o u7h�   h��jj��������@o�=@o u����  �@o�     �8o�M��}� u-3�u!h��j h�   h��j��������u̃���r  �M�+M�Q�U�R�  ���E�}� ��   �E��8 ��   j�M�U���P��������}� ti�	�M���M�U�E��<� t�M�U��E�u��D����ց}����?s2h�   h��jj�M�Q�8oR�������E��}� t�E��8o��M�U��E���M�    �   �}� ��   �}� }�U��ډU�E��;E�|:�M�������?s,h�   h��j�U��Rj�8oP�������E��}� u����D  �M�U��E���M�U��D�    �E�     �M��8o�j�U�R��������E�     3���   �} ��   h  h��jj�M�Q��������P�:�����E�}� ��   j h!  h��h��h8��U�R�E�P�������P�M�Q������P�y������U�+U�U�U��E��  �M����M��U������#U�R�E�P�����u�E������}��u���� *   j�M�Q��������}� tj�U�R��������E�     �E�^��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�8o�E��	�M����M��U��: tK�EP�M��R�EP��������u/�M���E���=t�U���M���u�E�+8o���뤋E�+8o���؋�]����������������������������������̋�U����E�    �E�E�} u3���   �M��E���E��t�M����M���h�  h��jj�U���R�5�����E��E��E��}� u
j	�T�����M�M�U�: ��   �E�Q��������E�h�  h��jj�U�R��
�����M���U��: t7j h�  h��h�h���E�Q�U�R�E��Q�����P�#������U���U�E����E��k����M��    �E���]��������������������������������������������������������������������������������̋�U���0�EP�M������3Ƀ} ���M�}� uh��j j:h@�j��������u̃}� u=�2���    j j:h@�h$�h��� �����E�    �M������E���   �M�������@�x u#�MQ�UR�U�����E��M�����E���   �	�E���E�Mf�f�U��E���t|�M��~����H�U��D��tS�M���M�U���u�E�    �M��?���E��j�M����U��9Mu�M���M؍M�����E��@��U�9Uu��h����E�9Eu�M�MԍM���
���E���E�    �M���
���EЋ�]���������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�N����]�������̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[������������������������������������������������������%X��%\��%`��%d��%h��%l��%p��%t��%x��%|��%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%Ē�%Ȓ�%̒�%В�%Ԓ�%ؒ�%ܒ�%���%��%��%��%��%���%���%���% ��%��%��%��%��%��%��%��% ��%$��%(��%,��%0��%4��%8��%<��%@��%D��%H��%L��%P��%T��%X��%\��%`��%d��%h��%l��%p��%t��%x��%|��%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%ē�%ȓ�%̓�%Г�%ԓ�%ؓ�%ܓ�%���%��%��%��%��%���%���%���̍M�������������������������T$�B������3��
���J�3��
������!����������������������������̍��������������������T$�B������3��S
������������������������������������̍M��{���T$�B�����3��
���8��������������̍M��K���T$�B�����3���	���h��a������������̍M�����T$�B�����3��	������1������������̍�x����������x������   ��x��������������Í�������������������������P�z���YÍ�$����y�����D����n����T$�B��d���3��"	���������������������������������������������������̍����������D���������0���������X���������M�������h���������l��������������� ���������������������������������������+��������J�����(����X����@����M����d����������������������������������!������������T$�B������3�� ���J�3������(��v���������������������������������������������������������������������������������̍���������T$�B�����3��~�������������������������������̍�������������������T$�B������3��3���@��������������������������������̋M�������M��������M�� �'����T$�B��$���3���������[����������������������̍M�	���M�������M���	���T$�B�����3������������������������������̋M���K����T$�B��$���3��N��������������������������������̍M��'	���������	���������	���������	���������������������T$�B������3������J�3������$��P���������������������������̍���������,������   ��,�����M���ËT$�B�����3��o���������������������������������̍M��G���������<���T$�B������3��&���J�3�������������������������������̋M�������M��������M�� �����T$�B��$���3��������K����������������������̋M�����T$�B�����3��������������������̋M������T$�B��$���3��a�������������������̍M�}���� ������   �� �����M�_���ËT$�B������3������������������������������������̍M��������������������   �������M�����ËT$�B������3�����T��'����������������������������������̍M����� ������   �� �����M����ËT$�B�����3��B������������������������������������̍M�M���T$�B�����3��������������������̋T$�B�����3������ ��Y��������������������̍M�������������   �������M����ËT$�B�����3�����\�������������������������������̋T$�B�����3��I���������������������������̍���������T$�B������3��������������������������������̋M������T$�B��$���3���������Q������������̋M�������T$�B��$���3��������!������������̋M������T$�B�����3��q�������������������̋M�����T$�B��$���3��A������������������̋M��d���T$�B��$���3�����H��������������̋M������T$�B��$���3��� ���x��a������������̋T$�B�����3�� ������9��������������������̍���������M��s����T$�B������3��v ���J�3��l ���L �������������������������̍M��G���������<���������1���M��)��������������������������������������������������@���������p�����������������������������X����������������������������������� ����������������0����y����H����n����l����c���������X���������M���������B���������7���������,��������!����,��������D��������\���� �������������������������������������������T$�B��4���3������J�3������x �4���������������������������������������������������������������������������������������������������������������̍M��7���������,���T$�B������3������J�3�������������������������������̍M������������`����������� ���T$�B������3������J�3������(�1����������������������������̍������ ���������y �������������������c ���������X ��������M ����H����B ����0����7 ����`����, ����x����! ��������� ���T$�B��@���3�� ����J�3�������T�v�������������������������������������������������̍MH������t���������P���������@�������������������,����������l����u�����T����j����������_����������T�������������������P�g���YË�$����0�����<����%����T$�B������3������J�3������������������������������������������������������������������������̍�P�������������������h����������������������������������}���������r�����L����g����������\���������Q�����4����F�����d����;�����|����0����������%���������������������������������������������H����������x���������� ����������0����������`���������������������������������������������������������������������D����u�����t����j����������_����������T�����,����I�����\����>����������3����������(���������������������������������4����������L����������d����������|���������T$�B������3���������E������������������������������������������������������������������������������������������������������������������������������������������������̍M��'������������������������T$�B������3�������J�3�������D�q����������������������������̍M������M��������t���������P���������,������������������������������������������������� �������������������t����Q�����P����t����������i����������0����������%����������������������������������(����������L���������p�����������������������������������������T$�B������3������J�3������p�"���������������������������������������������������������������������������������������������̍M,�7����M�/����M�'����M������M������M�������|���������d����������L����������4�������������������������������������������������������������$���������t���������D����M���T$�B������3��u����J�3��k����t������������������������������������������������������������������������̋M������T$�B��$���3������L�������������̋M�������T$�B��$���3�������|�Q������������̍M�������������   ��������M����ËT$�B������3�������������������������������������̍M�W������������   ��������M����ÍM������T$�B������3������J�3�����������������������������������̍M������T$�B������3�������,�Q������������̋M������M��@�����M���   �����M���   ��������������������z����T$�B������3��d����T���������������������������������̋M������M��@�����M���   �����M���   �����T$�B��$���3���������z���������������������̍M������T$�B������3�������	�A������������̍M�����M�����M�������M��(�����T$�B�����3��s����L	��������������������������������̋M���D����M��(�9����T$�B��$���3��#�����	�������������������������������̍M������T$�B�����3��������	�a������������̋M������M���_����T$�B��$���3�������	�&�����������������̋M��^����M�������M�� �K����T$�B�����3��[����8
������������������������̍M��|����������q����� ������   �� �����������P���Ë� ������   �� �����M�1���ËT$�B������3��������
�U��������������������������������̍����������T$�B�����3�������
��������������������������̍M�����M���������������������������������   ��������M����Í�d����d�����x���������������N����������C����T$�B������3��������
�h���������������������������������������������������̋M������T$�B��$���3������`�������������̋M��:����T$�B��$���3��a�������������������̍M����������������������v����������k����T$�B������3�����������������������������������̋M�������T$�B�����3��������Q������������̍M�g����� ������   �� �����M�����ËT$�B������3������D������������������������������̍M�����������������������   �������M�s���ËT$�B������3������������������������������������������̍M�����M���������������M��|����������q����� ����f����T$�B������3�������� ���������������������������̋M��:����T$�B�����3��a������������������̍M������� ������   �� �����M�n���ËT$�B�����3������P������������������������������̍M�����T$�B�����3���������Q������������̍M$�g����M�_����M�W����M��O����������D����������9����������.����������#����T$�B������3��]�����������������������������������������������̋T$�B�����3������P���������������������̍M��<����������I���������������������3���������(����T$�B��|���3������|�5��������������������������������̋M������T$�B��$���3��q�������������������̍M�������������   �������M�����ËT$�B�����3��"����������������������������������̍M�����M������ ������   �� ��������������Ë� ������   �� ���������������Ë� ������   �� �����M�����Í� ���������T$�B������3��k����D��������������������������������������������������������̋T$�B�����3����������������������������̍�����w����T$�B������3��������^�������������������������̍M�����T$�B�����3������8�!������������̍M�o����M�g����M�������M���������������   ��������M����ËT$�B������3��:����`��������������������������������������̍���������T$�B������3���������n�������������������������̍M������ ������   �� �����M����ËT$�B�����3�������������������������������������̍M�O����M������M������T$�B������3��A����@������������������������������̋M������T$�B��$���3��������������������̍M �����M�����M����������|���������q����T$�B������3�������+����������������������̋E�P�� ���Q�A�����ËT$�B�����3��e����`������������������̍M ������M������M�����������������M�������M�������T$�B������3�����������������������������������������̋T$�B�� ���3�������T�I��������������������̍M�W����M�O����� ����D����T$�B������3��~��������������������������������̋E�P�� ���Q������ËT$�B�����3��5����������������������̍M������T$�B��0���3��������������������̋T$�B�� ���3�������X�Y��������������������̍�������������������������������������������������T$�B������3��r������������������������������������̍M�G����T$�B�����3��1������������������̍M�������h��������������F�����d����y����������0������������������������������������������������ ����7����T$�B�����3������J�3������������������������������������������������������̍M�W����������L����������A����������6����� ����+��������� ��������������������
���������������� ����������P���������������������8����������h������������������������������������������������������������X���������p����{����������p����������e����������Z����������O����������D���������9�����$����.����T$�B��P���3�����������������������������������������������������������������������������������������������������������̍M����������������������������������������{�����$����p�����|����e����������Z����������O���������D����������9����������.����������#�����$���������<���������T���������l���������������������������������������������������������������� ���������D���������\���������t������������������������~����������s����T$�B��D���3��]�����������������������������������������������������������������������������������������������̍��������������������������������������������T$�B��,���3��������=������������������������̍����������L���������4����~�����d����s����������h����������]����������R����������G���������<�����<����1�����l����&�����$���������T��������������������������������������������������������������T$�B������3��������C��������������������������������������������������������������̍������t���������i�����4����^����������S���������H�����L����=�����d����2�����|����'����������������������������������� ����������0����������`�������������������������������H����������x���������������������������������������������������������������w����T$�B��`���3��a�����������������������������������������������������������������������������������̍�����������������������������������������������������4����������L����������d���������|���������������������������������������$��������������u���������j�����<����_�����T����T�����l����I����������>����������3����T$�B��H���3��������������������������������������������������������������������������������̍���������������������� ��������������������������������������0���������H����w���������l�����H����a�����x����V����������K����������@���������5�����0����*�����`������������������������	���������������� ����������8����������P����������h�������������������������������������������������������������������������������������z���������o�����4����d�����d����Y����������N����������C����������8�����$����-����������"��������������L���������|�����������������������������������������<����������T����������l����������������������������������������������������������������}���������r�����,����g�����D����\�����\����Q�����t����F����������;����������0����������%�����(����������������������������@����������X����������p���������T$�B������3���������M��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̍��������������������������������� ����������D����������t�����������������������������\����������������������������������{���������p���������e�����4����Z�����L����O�����p����D����������9����������.����� ����#�����0��������������������������������������������������H����������`����������x��������������������������������������������������T$�B��\���3������8�	����������������������������������������������������������������������������������������������������̍����������������	�������������������������������������(����������@����������X����������p������������������������������������������������<��������������z����������o�����$����d�����T����Y�����l����N����������C����������8����������-����������"��������������T$�B��<���3������|�����������������������������������������������������������������������������̍M�����������������������������������M��~�����H����s����������h�����@����]�����$����9�����X����G����������<����������1�����0����&��������������H���������x���������������������������������������������������������������D����������t�������������������,���������\����������������������������������v����������k����������`���������U�����@����J�����p����?����������4�����(����)�����X��������������������������������������������������� ��������������������<����������l����������T����������������������������������������������������������� ����y���������鳿����P���������x���靿���������M����������B����������7����� ����,�����$����!�����`���������H���������x���� ���������������������m�����0��������������������T��������������������l������������������T$�B��0���3������J�3������x��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̍M��*����T$�B�J�3������"����������������̍M�������T$�B�J�3��d����\"�����������������̍M��ʻ���T$�B�J�3��4�����"����������������̋T$�B�J�3�������'������������������������̍M�������T$�B�J�3��������,�T���������������̡4v����4vËT$�B�J�3������0.��������������������������̍M��[����T$�B�J�3��d�����/�����������������̍M��+����T$�B�J�3��4����00����������������̍M�������T$�B�J�3������`1����������������̍M�������T$�B�J�3��������1�T��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �����󫹔c�<���h��������_^[���   ;�������]������������������������U����   SVW��@����0   ������j ��c�����_^[���   ;��Ʃ����]������������������̋�U���h����h�������]������������������̋�U��Q3��E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �����󫹔c�j���_^[���   ;��(�����]��������������������̋�U���h�}���]���������������̋�U��i�؈��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           p�                                                                                                                                                                                                                                                                �� ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            I�Ռ,�W��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            F�	�                                                                                                                                                                                                                                                                    ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    6ڀL       s   t� te bad allocation                           ?                             @   �                       0   @   �  �      0                                 @   �                 LOD-Object          I T E R A T O R   L I S T   C O R R U P T E D !             c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   9 . 0 \ v c \ i n c l u d e \ x u t i l i t y                                   �? @F     ���R���u���� �ɢE�1�ҙS�}�֤~�ݓ������O�����a����������ϡ՛                            level [      ]
  ,  range [     
       center      DEF      LOD{
  c:\program files (x86)\cinema 4d r10\plugins\vrmlexporter\source\object\lod.cpp                 }
  ]
  lod.tif     Olevelofdetail      VRMLExporter-LOD        c:\program files (x86)\cinema 4d r10\plugins\vrmlexporter\source\object\lod.h                   0���V���u���g� �ɢE�1�ҙS�h���~�6������O�����a���������ϡ՛                                H�q�V���u���g� �ɢE�1�ҙS�h���~�6�                    c:\program files (x86)\microsoft visual studio 9.0\vc\include\xdebug                `�:�ɧ        l i s t   e r a s e   i t e r a t o r   o u t s i d e   r a n g e                       c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   9 . 0 \ v c \ i n c l u d e \ l i s t                             l i s t   i n s e r t   i t e r a t o r   o u t s i d e   r a n g e                 " o u t   o f   r a n g e "         s t d : : l i s t < c l a s s   L O D m g m t   * , c l a s s   s t d : : a l l o c a t o r < c l a s s   L O D m g m t   * >   > : : _ C o n s t _ i t e r a t o r < 1 > : : o p e r a t o r   *                                               ( " S t a n d a r d   C + +   L i b r a r i e s   O u t   o f   R a n g e " ,   0 )                     l i s t   i t e r a t o r   n o t   d e r e f e r e n c a b l e                 s t d : : l i s t < c l a s s   L O D m g m t   * , c l a s s   s t d : : a l l o c a t o r < c l a s s   L O D m g m t   * >   > : : _ C o n s t _ i t e r a t o r < 1 > : : o p e r a t o r   + +                                             l i s t   i t e r a t o r   n o t   i n c r e m e n t a b l e                   s t d : : l i s t < c l a s s   L O D m g m t   * , c l a s s   s t d : : a l l o c a t o r < c l a s s   L O D m g m t   * >   > : : _ C o n s t _ i t e r a t o r < 1 > : : o p e r a t o r   - -                                             l i s t   i t e r a t o r   n o t   d e c r e m e n t a b l e               " i n v a l i d   a r g u m e n t "                 s t d : : l i s t < c l a s s   L O D m g m t   * , c l a s s   s t d : : a l l o c a t o r < c l a s s   L O D m g m t   * >   > : : _ C o n s t _ i t e r a t o r < 1 > : : _ C o m p a t                                             ( " S t a n d a r d   C + +   L i b r a r i e s   I n v a l i d   A r g u m e n t " ,   0 )                     l i s t   i t e r a t o r s   i n c o m p a t i b l e               list<T> too long    ���0�    ��t�0�    ����    c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   9 . 0 \ v c \ i n c l u d e \ x s t r i n g                               i n v a l i d   n u l l   p o i n t e r             �zBH�Q@���?���?  �  ��  @�   �   A  @@NavigationInfo-Object       visibilityLimit     type ["     "]
 speed   headlight       avatarSize [    ,   NavigationInfo{ 
       NONE    FLY EXAMINE     WALK    ANY FALSE   TRUE        ����K���u����� �ɢE�1�ҙS�h���~�6������O�����a�W��������ϡ՛                            navinfo.tif     onavigationinfo     VRMLExporter-NavigationInfo             c:\program files (x86)\cinema 4d r10\plugins\vrmlexporter\source\object\navigationinfo.h                    ������)�K���)�j�k�        

  #   Date:   # CINEMA4D File:        ## Produced by Florian's VRML Plugin, Version alpha_0.2 
               #VRML V2.0 utf8

       -   children [
     rotation    scale   translation      Transform { 
             @              �?        -DT�!	@              �                    fvrmlexport     wrl VRML Exporter   c:\program files (x86)\cinema 4d r10\plugins\vrmlexporter\source\scenesaver\vrmlexp.h                    �\�V���u���g� �ɢE�1�ҙS�h���~�6���                ���V���u���g� �ɢE�1�ҙS�h���~�6�,�                #Couldn't find/copy Textur:         \tex\   \maps\  \   /   �����@�)�K�5�)�j�k�            c:\program files (x86)\cinema 4d r10\plugins\vrmlexporter\source\scenesaver\vrmlexp.cpp                       �@l i s t   s p l i c e   i t e r a t o r   o u t s i d e   r a n g e                 ( " _ P o s   <   s i z e ( ) " ,   0 )             s t d : : v e c t o r < c l a s s   s t d : : l i s t < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   > , c l a s s   s t d : : a l l o c a t o r < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   >   >   > : : _ I t e r a t o r < 1 > , c l a s s   s t d : : a l l o c a t o r < c l a s s   s t d : : l i s t < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   > , c l a s s   s t d : : a l l o c a t o r < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   >   >   > : : _ I t e r a t o r < 1 >   >   > : : o p e r a t o r   [ ]                                                                                                                                                                                                               v e c t o r   s u b s c r i p t   o u t   o f   r a n g e                   c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   9 . 0 \ v c \ i n c l u d e \ v e c t o r                                 s t d : : l i s t < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   > , c l a s s   s t d : : a l l o c a t o r < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   >   >   > : : _ C o n s t _ i t e r a t o r < 1 > : : _ C o m p a t                                                                                                   s t d : : l i s t < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   > , c l a s s   s t d : : a l l o c a t o r < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   >   >   > : : _ C o n s t _ i t e r a t o r < 1 > : : o p e r a t o r   *                                                                                                     s t d : : l i s t < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   > , c l a s s   s t d : : a l l o c a t o r < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   >   >   > : : _ C o n s t _ i t e r a t o r < 1 > : : o p e r a t o r   + +                                                                                                           s t d : : l i s t < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   > , c l a s s   s t d : : a l l o c a t o r < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   >   >   > : : _ C o n s t _ i t e r a t o r < 1 > : : o p e r a t o r   - -                                                                                                           v e c t o r   e r a s e   i t e r a t o r   o u t s i d e   r a n g e                   vector<T> too long      v e c t o r   i n s e r t   i t e r a t o r   o u t s i d e   r a n g e                 s t d : : _ V e c t o r _ c o n s t _ i t e r a t o r < c l a s s   s t d : : l i s t < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   > , c l a s s   s t d : : a l l o c a t o r < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   >   >   > : : _ I t e r a t o r < 1 > , c l a s s   s t d : : a l l o c a t o r < c l a s s   s t d : : l i s t < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   > , c l a s s   s t d : : a l l o c a t o r < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   >   >   > : : _ I t e r a t o r < 1 >   >   > : : _ V e c t o r _ c o n s t _ i t e r a t o r                                                                                                                                                                                                                             ( " _ P v e c t o r   = =   N U L L   | |   ( ( ( _ M y v e c   * ) _ P v e c t o r ) - > _ M y f i r s t   < =   _ P t r   & &   _ P t r   < =   ( ( _ M y v e c   * ) _ P v e c t o r ) - > _ M y l a s t ) " ,   0 )                                                 s t d : : _ V e c t o r _ c o n s t _ i t e r a t o r < c l a s s   s t d : : l i s t < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   > , c l a s s   s t d : : a l l o c a t o r < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   >   >   > : : _ I t e r a t o r < 1 > , c l a s s   s t d : : a l l o c a t o r < c l a s s   s t d : : l i s t < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   > , c l a s s   s t d : : a l l o c a t o r < c l a s s   s t d : : b a s i c _ s t r i n g < c h a r , s t r u c t   s t d : : c h a r _ t r a i t s < c h a r > , c l a s s   s t d : : a l l o c a t o r < c h a r >   >   >   > : : _ I t e r a t o r < 1 >   >   > : : _ C o m p a t                                                                                                                                                                                                                       v e c t o r   i t e r a t o r s   i n c o m p a t i b l e               i n v a l i d   i t e r a t o r   r a n g e                 c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   9 . 0 \ v c \ i n c l u d e \ m e m o r y                                 Do you want to replace the older file:           with the new one?      Dataconflict!     �B�������^��L>���=ROUTE   -POS-INTERP.value_changed TO        .set_translation

      ROUTE Timer.fraction_changed TO         -POS-INTERP.set_fraction
       ] } 
   Position . Z    Position . Y    Position . X    keyValue [ 
    ] 
 ,   key[ 
  -POS-INTERP PositionInterpolator { 
          zD      �?             @�@    �_c�  4&�k�    �_cX  4&�kC    -ROT-INTERP.value_changed TO        .set_rotation

     -ROT-INTERP.set_fraction
       ] }

       ����MbP?    
] 
    key [ 
     -ROT-INTERP OrientationInterpolator {
          }

       loop TRUE
          cycleInterval               stopTime 0
             startTime 0
      DEF Timer TimeSensor {
     # Camera, hier noch als Bsp. noch nicht implementiert 
             point [     coord DEF       -COORD Coordinate { 
       solid FALSE
    geometry DEF    -GEOMETRY IndexedFaceSet {
         , -1,
  coordIndex  [ 
     vector[     normal Normal {
    normalPerVertex TRUE 
      texCoord     USE    -TEXCOORD1
     ,
    ��point [ 
   texCoord DEF    -TEXCOORD    TextureCoordinate { 
      , -1,
      texCoordIndex    [ 
    texCoordIndex [ 
       normalIndex [ 
     material Material { }
      appearance Appearance {
        appearance  USE     " }
    texture DEF TEXTURE_         ImageTexture{ url "maps/       texture USE TEXTURE_        } 
 transparency    shininess       specularColor       diffuseColor    ambientIntensity         
  material Material { 
       appearance  DEF      Appearance {
      )\���(�?        �z�G��?        333333�?              $@           ����?           `ff�?    -SHAPE Shape {
     c:\program files (x86)\cinema 4d r10\resource\_api\c4d_resource.cpp                 #   M_EDITOR        c:\program files (x86)\cinema 4d r10\resource\_api\c4d_baseobject.cpp               $���    ��,�    �����         �8�9�C    res 0�;�        c:\program files (x86)\cinema 4d r10\resource\_api\c4d_string.cpp                B   KB  MB           �@     GB    %s  c:\program files (x86)\cinema 4d r10\resource\_api\c4d_file.cpp             H� �1�@�)�K�5�)�j���                 �f@              Y@    `���1�@�)�K�5�)�j�k�        x�v� ��f�ߪ8�����9���P�            ��~�1�@�)�K�5�)�j�ܞ        ~       ,��1�@�)�K�5�)�j��ڪħ}�p�����7���`���;��                         �Ngm��C              �A    ���� ����ߪ8�{���9�����            c:\program files (x86)\cinema 4d r10\resource\_api\c4d_customdatatype.cpp               ��׏,�c��9�����֩        c:\program files (x86)\cinema 4d r10\resource\_api\c4d_libs\lib_ngon.cpp                   ?    c:\program files (x86)\cinema 4d r10\resource\_api\c4d_pmain.cpp                unknown     exception:         f:\dd\vctools\crt_bld\self_x86\crt\src\xdebug           string too long     invalid string position     D���0�    invalid string argument     ����0�        f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ x s t r i n g                                     ��7�7�    �U�    csm�               �                \��ɧ    Unknown exception       t���ɧ    ��]�ɧ    ,���ɧ    . . .       A s s e r t i o n   F a i l e d         E r r o r       W a r n i n g       �Z�Z\Z    f:\dd\vctools\crt_bld\self_x86\crt\src\dbgrpt.c                 ( " T h e   h o o k   f u n c t i o n   i s   n o t   i n   t h e   l i s t ! " , 0 )                       p f n N e w H o o k   ! =   N U L L             _ C r t S e t R e p o r t H o o k W 2               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g r p t . c                           m o d e   = =   _ C R T _ R P T H O O K _ I N S T A L L   | |   m o d e   = =   _ C R T _ R P T H O O K _ R E M O V E                           M i c r o s o f t   V i s u a l   C + +   D e b u g   L i b r a r y                     _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r                     w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                   ( * _ e r r n o ( ) )           D e b u g   % s ! 
 
 P r o g r a m :   % s % s % s % s % s % s % s % s % s % s % s % s 
 
 ( P r e s s   R e t r y   t o   d e b u g   t h e   a p p l i c a t i o n )                                     
 M o d u l e :         
 F i l e :         
 L i n e :         
 
     E x p r e s s i o n :               
 
 F o r   i n f o r m a t i o n   o n   h o w   y o u r   p r o g r a m   c a n   c a u s e   a n   a s s e r t i o n 
 f a i l u r e ,   s e e   t h e   V i s u a l   C + +   d o c u m e n t a t i o n   o n   a s s e r t s .                                                     m e m c p y _ s ( s z S h o r t P r o g N a m e ,   s i z e o f ( T C H A R )   *   ( 2 6 0   -   ( s z S h o r t P r o g N a m e   -   s z E x e N a m e ) ) ,   d o t d o t d o t ,   s i z e o f ( T C H A R )   *   3 )                                                 < p r o g r a m   n a m e   u n k n o w n >                 w c s c p y _ s ( s z E x e N a m e ,   2 6 0 ,   L " < p r o g r a m   n a m e   u n k n o w n > " )                       _ _ c r t M e s s a g e W i n d o w W           s i z e I n B y t e s   > =   c o u n t             s r c   ! =   N U L L       m e m c p y _ s             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m e m c p y _ s . c                       d s t   ! =   N U L L       m e m m o v e _ s           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m e m m o v e _ s . c                         (   t i m p   ! =   N U L L   )         _ c t i m e 6 4 _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c t i m e 6 4 . c                         (   (   b u f f e r   ! =   N U L L   )   & &   (   s i z e I n C h a r s   >   0   )   )                       _ c t i m e 6 4         ( " I n v a l i d   f i l e   d e s c r i p t o r .   F i l e   p o s s i b l y   c l o s e d   b y   a   d i f f e r e n t   t h r e a d " , 0 )                                   ( _ o s f i l e ( f h )   &   F O P E N )           _ c l o s e     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c l o s e . c                     ( f h   > =   0   & &   ( u n s i g n e d ) f h   <   ( u n s i g n e d ) _ n h a n d l e )                     ( _ o s f i l e ( f i l d e s )   &   F O P E N )               ( f i l d e s   > =   0   & &   ( u n s i g n e d ) f i l d e s   <   ( u n s i g n e d ) _ n h a n d l e )                         _ f s t a t 6 4 i 3 2       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f s t a t 6 4 . c                         ( b u f   ! =   N U L L )               s t r c p y _ s ( p f d - > n a m e ,   ( s i z e o f ( p f d - > n a m e )   /   s i z e o f ( p f d - > n a m e [ 0 ] ) ) ,   w f d . c F i l e N a m e )                                     ( s z W i l d   ! =   N U L L )         ( s i z e o f ( p f d - > n a m e )   < =   s i z e o f ( w f d . c F i l e N a m e ) )                     _ f i n d f i r s t 6 4 i 3 2               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f i n d f 6 4 . c                         ( p f d   ! =   N U L L )           _ f i n d n e x t 6 4 i 3 2         ( ( H A N D L E ) h F i l e   ! =   I N V A L I D _ H A N D L E _ V A L U E )                         �?      �?3      3            �      0C       �       ��                                  f:\dd\vctools\crt_bld\self_x86\crt\src\dllcrt0.c            f:\dd\vctools\crt_bld\self_x86\crt\src\onexit.c             ( s t r i n g   ! =   N U L L )         _ v s p r i n t f _ l       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v s p r i n t f . c                       ( f o r m a t   ! =   N U L L )         _ v s c p r i n t f _ h e l p e r               (   ( _ S t r e a m - > _ f l a g   &   _ I O S T R G )   | |   (   f n   =   _ f i l e n o ( _ S t r e a m ) ,   (   ( _ t e x t m o d e _ s a f e ( f n )   = =   _ _ I O I N F O _ T M _ A N S I )   & &   ! _ t m _ u n i c o d e _ s a f e ( f n ) ) ) )                                                       ( s t r e a m   ! =   N U L L )         f p u t s           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f p u t s . c                     f:\dd\vctools\crt_bld\self_x86\crt\src\_file.c          Client  Ignore  CRT Normal  Free    �o�o�o�o�o    Error: memory allocation: bad memory block type.
           Invalid allocation size: %Iu bytes.
        Client hook allocation failure.
        Client hook allocation failure at file %hs line %d.
                f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g h e a p . c                         _ C r t C h e c k M e m o r y ( )           _ c a l l o c _ d b g _ i m p l         ( _ H E A P _ M A X R E Q   /   n N u m )   > =   n S i z e                 _ p F i r s t B l o c k   = =   p O l d B l o c k               _ p L a s t B l o c k   = =   p O l d B l o c k                 f R e a l l o c   | |   ( ! f R e a l l o c   & &   p N e w B l o c k   = =   p O l d B l o c k )                       Error: possible heap corruption at or near 0x%p                 p O l d B l o c k - > n L i n e   = =   I G N O R E _ L I N E   & &   p O l d B l o c k - > l R e q u e s t   = =   I G N O R E _ R E Q                                 _ C r t I s V a l i d H e a p P o i n t e r ( p U s e r D a t a )                       The Block at 0x%p was allocated by aligned routines, use _aligned_realloc()                     Error: memory allocation: bad memory block type.

Memory allocated at %hs(%d).
                 Invalid allocation size: %Iu bytes.

Memory allocated at %hs(%d).
              Client hook re-allocation failure.
         Client hook re-allocation failure at file %hs line %d.
             _ r e c a l l o c _ d b g           ( _ H E A P _ M A X R E Q   /   c o u n t )   > =   s i z e                 _ e x p a n d _ d b g       p U s e r D a t a   ! =   N U L L           _ p F i r s t B l o c k   = =   p H e a d           _ p L a s t B l o c k   = =   p H e a d             p H e a d - > n B l o c k U s e   = =   n B l o c k U s e               p H e a d - > n L i n e   = =   I G N O R E _ L I N E   & &   p H e a d - > l R e q u e s t   = =   I G N O R E _ R E Q                                 HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.
                           HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.

Memory allocated at %hs(%d).
                                     HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.
                               HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.

Memory allocated at %hs(%d).
                                         _ B L O C K _ T Y P E _ I S _ V A L I D ( p H e a d - > n B l o c k U s e )                     Client hook free failure.
      The Block at 0x%p was allocated by aligned routines, use _aligned_free()                _ m s i z e _ d b g         %hs located at 0x%p is %Iu bytes long.
             %hs located at 0x%p is %Iu bytes long.

Memory allocated at %hs(%d).
                   HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.
                               HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.

Memory allocated at %hs(%d).
                                 DAMAGED     _heapchk fails with unknown return value!
          _heapchk fails with _HEAPBADPTR.
       _heapchk fails with _HEAPBADEND.
       _heapchk fails with _HEAPBADNODE.
          _heapchk fails with _HEAPBADBEGIN.
         _ C r t S e t D b g F l a g             ( f N e w B i t s = = _ C R T D B G _ R E P O R T _ F L A G )   | |   ( ( f N e w B i t s   &   0 x 0 f f f f   &   ~ ( _ C R T D B G _ A L L O C _ M E M _ D F   |   _ C R T D B G _ D E L A Y _ F R E E _ M E M _ D F   |   _ C R T D B G _ C H E C K _ A L W A Y S _ D F   |   _ C R T D B G _ C H E C K _ C R T _ D F   |   _ C R T D B G _ L E A K _ C H E C K _ D F )   )   = =   0 )                                                                                 _ C r t D o F o r A l l C l i e n t O b j e c t s               p f n   ! =   N U L L       Bad memory block found at 0x%p.
        Bad memory block found at 0x%p.

Memory allocated at %hs(%d).
              _ C r t M e m C h e c k p o i n t           s t a t e   ! =   N U L L           n e w S t a t e   ! =   N U L L         o l d S t a t e   ! =   N U L L         _ C r t M e m D i f f e r e n c e           Object dump complete.
      crt block at 0x%p, subtype %x, %Iu bytes long.
             normal block at 0x%p, %Iu bytes long.
          client block at 0x%p, subtype %x, %Iu bytes long.
              {%ld}   %hs(%d) :       #File Error#(%d) :      Dumping objects ->
      Data: <%s> %s
     _ p r i n t M e m B l o c k D a t a             %.2X    Detected memory leaks!
     Total allocations: %Id bytes.
          Largest number used: %Id bytes.
        %Id bytes in %Id %hs Blocks.
       _ C r t M e m D u m p S t a t i s t i c s           o f f s e t   = =   0   | |   o f f s e t   <   s i z e                 _ a l i g n e d _ o f f s e t _ m a l l o c _ d b g             I S _ 2 _ P O W _ N ( a l i g n )           _ a l i g n e d _ o f f s e t _ r e a l l o c _ d b g               Damage before 0x%p which was allocated by aligned routine
              The block at 0x%p was not allocated by _aligned routines, use realloc()                 _ a l i g n e d _ o f f s e t _ r e c a l l o c _ d b g                 The block at 0x%p was not allocated by _aligned routines, use free()                _ a l i g n e d _ m s i z e _ d b g             m e m b l o c k   ! =   N U L L         Unknown Runtime Check Error
       Stack memory around _alloca was corrupted
         A local variable was used before it was initialized
           Stack memory was corrupted
        A cast to a smaller data type has caused a loss of data.  If this was intentional, you should mask the source of the cast with the appropriate bitmask.  For example:  
	char c = (i & 0xFF);
Changing the code in this way will not affect the quality of the resulting optimized code.
                                                            The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.
                                                `�����p�L�                   Stack around the variable ' ' was corrupted.    The variable '  ' is being used without being initialized.                                  Run-Time Check Failure #%d - %s         Unknown Module Name     Unknown Filename        R u n - T i m e   C h e c k   F a i l u r e   # % d   -   % s                   R u n t i m e   C h e c k   E r r o r . 
    U n a b l e   t o   d i s p l a y   R T C   M e s s a g e .                           Stack corrupted near unknown variable               Stack area around _alloca memory reserved by this function is corrupted
                %s%s%s%s    >   %s%s%p%s%ld%s%d%s       Stack area around _alloca memory reserved by this function is corrupted                 
Address: 0x    
Size:      
Allocation number within this function:            
Data: <    wsprintfA   user32.dll      A variable is being used without being initialized.             Stack around _alloca corrupted          Local variable used before initialization           Stack memory corruption     Cast to smaller type causing loss of data           Stack pointer corruption        č��t�@��    f:\dd\vctools\crt_bld\self_x86\crt\prebuild\misc\i386\chkesp.c              The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.                                              ��bad exception   ��
�ɧ    EncodePointer   K E R N E L 3 2 . D L L         DecodePointer   f:\dd\vctools\crt_bld\self_x86\crt\src\tidtable.c           FlsFree     FlsSetValue     FlsGetValue     FlsAlloc    �i j        _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   0 x 0 0 0 1 0 0 0 0 ,   0 x 0 0 0 3 0 0 0 0 )                       _ s e t d e f a u l t p r e c i s i o n                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n t e l \ f p 8 . c                                �~PA           ���GA    IsProcessorFeaturePresent       KERNEL32    s i z e I n B y t e s   >   0           _ c f t o e _ l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ c v t . c                         b u f   ! =   N U L L       e+000   s t r c p y _ s ( p ,   ( s i z e I n B y t e s   = =   ( s i z e _ t ) - 1   ?   s i z e I n B y t e s   :   s i z e I n B y t e s   -   ( p   -   b u f ) ) ,   " e + 0 0 0 " )                                       s i z e I n B y t e s   >   ( s i z e _ t ) ( 3   +   ( n d e c   >   0   ?   n d e c   :   0 )   +   5   +   1 )                           _ c f t o e 2 _ l           s i z e I n B y t e s   >   ( s i z e _ t ) ( 1   +   4   +   n d e c   +   6 )                     _ c f t o a _ l         _ c f t o f _ l         _ c f t o f 2 _ l       _ c f t o g _ l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ e h \ t y p n a m e . c p p                             p N o d e - > n e x t   ! =   N U L L           s t r c p y _ s   ( ( c h a r   * ) ( ( t y p e _ i n f o   * ) _ T h i s ) - > _ m _ d a t a ,   l e n + 2 ,   ( c h a r   * ) p T m p U n d N a m e )                                 t y p e _ i n f o : : _ N a m e _ b a s e               s t r c p y _ s   ( p T m p T y p e N a m e ,   l e n + 2 ,   ( c h a r   * ) p T m p U n d N a m e )                       t y p e _ i n f o : : _ N a m e _ b a s e _ i n t e r n a l                 ( L " B u f f e r   i s   t o o   s m a l l "   & &   0 )               B u f f e r   i s   t o o   s m a l l           ( ( ( _ S r c ) ) )   ! =   N U L L             s t r c p y _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s c p y _ s . i n l                           ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n B y t e s ) )   >   0                     f:\dd\vctools\crt_bld\self_x86\crt\src\mlock.c              f M o d e   = =   _ C R T D B G _ R E P O R T _ M O D E   | |   ( f M o d e   &   ~ ( _ C R T D B G _ M O D E _ F I L E   |   _ C R T D B G _ M O D E _ D E B U G   |   _ C R T D B G _ M O D E _ W N D W ) )   = =   0                                                 _ C r t S e t R e p o r t M o d e               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g r p t t . c                         n R p t T y p e   > =   0   & &   n R p t T y p e   <   _ C R T _ E R R C N T                   _ C r t S e t R e p o r t F i l e               _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g                             w c s c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )                                         e   =   m b s t o w c s _ s ( & r e t ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                               s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )                           s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                 %s(%d) : %s         s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ n " )                          s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ r " )                   s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )                         s t r c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   " A s s e r t i o n   f a i l e d :   "   :   " A s s e r t i o n   f a i l e d ! " )                                     Assertion failed!       Assertion failed:       _CrtDbgReport: String too long or IO Error          s t r c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                   , Line      <file unknown>      Second Chance Assertion Failed: File            _ i t o a _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )                   _ V C r t D b g R e p o r t A           w c s t o m b s _ s ( & r e t ,   s z a O u t M e s s a g e ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                               _CrtDbgReport: String too long or Invalid characters in String                  s t r c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )                                           w c s t o m b s _ s ( ( ( v o i d   * ) 0 ) ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                                 w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )                       % s ( % d )   :   % s       w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ n " )                        w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ r " )                 w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )                         w c s c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   L " A s s e r t i o n   f a i l e d :   "   :   L " A s s e r t i o n   f a i l e d ! " )                                     A s s e r t i o n   f a i l e d !           A s s e r t i o n   f a i l e d :                   w c s c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                 
   ,   L i n e         < f i l e   u n k n o w n >             S e c o n d   C h a n c e   A s s e r t i o n   F a i l e d :   F i l e                         _ i t o w _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )                   _ V C r t D b g R e p o r t W           _ g e t _ e r r n o             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d o s m a p . c                       p V a l u e   ! =   N U L L         _ g e t _ d o s e r r n o           CorExitProcess      m s c o r e e . d l l       _ w p g m p t r   ! =   N U L L         _ g e t _ w p g m p t r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c r t 0 d a t . c                         _ p g m p t r   ! =   N U L L           _ g e t _ p g m p t r       s i g n a l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w i n s i g . c                       ( " I n v a l i d   s i g n a l   o r   e r r o r " ,   0 )                 f:\dd\vctools\crt_bld\self_x86\crt\src\winsig.c             r a i s e       GetProcessWindowStation     GetUserObjectInformationW       GetLastActivePopup      GetActiveWindow     MessageBoxW     U S E R 3 2 . D L L         _ s w p r i n t f       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s w p r i n t f . c                       w c s c p y _ s         ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n W o r d s ) )   >   0                               �?    ���?     ��?    �D�?    ��?     ��?    @��?    @W�?     �?    ���?    ���?    �w�?    �A�?    ��?    @��?    ���?    �q�?    �?�?     �?    @��?     ��?    �}�?    �N�?    @ �?    ���?    ���?     ��?     m�?    �A�?    ��?    ���?    ���?    ���?     q�?    �H�?     !�?    ���?     ��?    ���?     ��?    �a�?    �<�?     �?     ��?    @��?    @��?    @��?    �g�?    �E�?    @$�?     �?     ��?    ���?    @��?    ���?     b�?    �B�?     $�?    ��?    @��?    ���?     ��?    ���?     r�?    @U�?     9�?     �?    @�?     ��?    ���?    ���?    @��?     {�?    �`�?     G�?    �-�?     �?     ��?    @��?    ���?    @��?     ��?    @��?    �i�?     R�?     ;�?     $�?     �?    ���?    @��?     ��?     ��?    @��?    ���?    @s�?    @^�?    @I�?    @4�?    ��?    @�?     ��?     ��?     ��?    @��?    ���?    @��?     ��?     n�?     [�?    @H�?    �5�?    @#�?     �?     ��?     ��?    @��?    ���?     ��?    ���?    @��?    @��?    @s�?    @b�?    �Q�?     A�?    �0�?    @ �?     �?      �?                          �a���?���F��<=  z1%�?�Vd?E=  ��b�?�6��\�M=  ���?p�9t^�<= �\c�N�?	�ʽ��J= �3���?�/��N=  �b�?DZ.�0=  �Ohe�?�?���0=  ]3��?��`$= @�׹ƻ?X&eB�E= ���rr�?\�3#�.J= ��׌�?��C5= �3:���?Ltm��YE= @�'z+�?�"e���=  tLVv�?p��$��M= `�dH��?h6_~��(= `x��?��Y�O= ���YL�?wJ�Q�\C= ��jU��?�Vш4= �+0��?e���37.= `�2�?�⋱�K= `���I�?)-��W�0=  -�Ƀ�?���*D= ���D��?7Tf(��G= �6	�x�?Y��8= ��%��?�E�<= ��w��?�~�?= �Ґ�C�?]���u�<= P��W��?>#�4�<  ��Xq�?���B�J= �_D��?m��K��F= ��Ԛ�?��s7�E= @�[-�?K>�d�:= ��g��?Z}�=\uI= �s�~Q�?�g:"(�N= �'��?9�~$O1=  ��q�?�n�1��%= p)k� �?v�ʌ�= `�X:��?�q.W�� = Pi���?g���>�M= ��[��?ֲa
��M= �_�3�?֍,�uXO= `Ɏ/��?���1w<= �>'eH�?`�	J�J= x~��? �&= n�`Y�?��˖��C= 0����?�]��/= # �g�?u�P�= �����?���,l�C= �5��q�?ᕎ�	= @Dӳ��?�-[�@= pt�4z�? �فpnJ= ���l��?�i�.Eg�< �y~�?�?�O�^'= (T�t��?�
�x;�;=  �P��?�R�RF= ��&�?X��ɣN= �J��@�?��~��= Ht=c��?Az�U"= ��nB��?U_l�j7= ��]���?q���BD=  �h<�?z�)�t'= �Z�#z�?��0�L= @5��ڿS�OO�F� ��ڿ���ۓ�D� 0���ٿ��= �n�  �W9!ٿ?�j>� 0�"�ؿ�؍� �I� �Q�n0ؿ�Hn&�E� �:�׿E7D���5� ��7�A׿��%@� @���ֿ* ��Z+A� �S��Tֿ�rJ� �D� @ӑ��տ����NT?� �w3�kտr�1�9�  �]��ԿF�K�m�8� �C!`�Կ1y2�Y�� @��Կ*�(<j�  䃝ӿV�CD� p��,ӿ1���n� ��ҿ2�=l�7� 0���IҿO���	x*�  �l@�ѿ2��>�FE� �O�5iѿ���4�Q!� �?:	�п�C	 ��+� pڌX�п��xO,�C�  �"пA��ri<� �q~�_Ͽ�R� v=� �=	~�ο����o6� @m�P�Ϳ	 ���d+� �>��̿9Ȓ���� �[\�˿8�B��'� ����&˿�i�[J� ��Z�Oʿ�b�n�E� �D�E}ɿ�Ugc@� �H	��ȿUZ�d��L�  "� �ǿ=��Dj!�  ��ǿ��Vm�:A� @��`3ƿ�~%�3�  k��cſ�"�7M�  ����Ŀ��p��>� �)%��ÿ\�����B� ��jx�¿#6HQ;� `t�-¿=]P��H0� �;T�a�����ָE�  &�����a-#��K� �V\���Vb���4M� @������U@�  X�x�����55� @���캿D��=� �iI�^��Gי��'7� ��A�Է�U�����N�  ��<N���>Ҫ1� ���Gƴ��O\�C� @��+B���g:IB� @Z�u�������}M� ����:��(T��!1� ���n���]vQ<)8�  h׾o��$�|�f+� ����x��2S��74�  U".���mœFB*� �6�I���KS�_D�   �5��M�-�C�  z1}B����K� G�  �c��?�Of��F�  �L,��s�X4I+�  xm�	w�$��V�cE�                      �?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    �
�?    �
�?    @
�?     
�?    �	�?    �	�?    @	�?     	�?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    � �?    � �?    @ �?      �?                          �|)P!?Ua0�		!=   �+34?�2��Q	=  �`��??7;W��J=  `�7�E?��'a %C=  ��MkK?�*��b<=  0ɘP?*�,�z?=  d|S?�K�T'�K=   �R_V?�b���F=  p^�BY?�����E&=  �9&\?�߇�N9=  p��	_?߭Eb2]A=  ���`?��f#I=  ���hb?O2�H`3=  ����c?e2��a�1=  �ԆLe?2���RM=  ����f?A�3�_:=  @�0h?[��2ieO=  ����i?�1r�K=  ���k?����Σ-=  ���l?���̈[8=  �yQ�m?>�|W8A=  �՛ko?�>qݲN=  ���np?z m{M=  t�)(q?m,�S�D=   E`�q?��}e?=  ԩ��r?�}~:f�E=  P��Ss?����&�A=  ��&t?,&��8=  ��t�t?�eѴN�@=  PS�u?^p?o4�0=  �!9v?�W�?N=  <��v?+�#�GYM=  H�w?qC���@=  ��Pex?0&ے=  X��y?���8 =  <8�y?!({=�H=   ���z?�d,G�B=  ��6K{?ҝ��E	M=  �¾|?w�3�1�!=  ��L�|?��^X-F=  �<�w}?0��!�O=  ��y1~?|"į�Q<=  $�~?��k�f@=  �+��?��b�UC=  ��4/�?*�K_�<*=  <��t�?�̍xI=  2�р?wY�V%A+=  ���.�?x+s7�E=  8#o��?�e��fE=  �|R�?Ks޸�E=  T�8E�?�=��(=  ��!��?��)��G=  ���?#F؇K=  V�[�?��C�<  :︃?k�V���I=  ����?����YH=  ���r�?q��4';=  .~�τ?��=�S7=  �'�,�?7���X�#=  4�ԉ�?C��k��7=  bB��?��EpC=  B��C�?'�2xk==  蠆?̸WU�A=  xm�	w�$��V�cE�  ̑ʭv�K��[��7�  �G�Qv�e$�l�F�  ����u��y�ԏ�H�  �gԙu�|��ǣ%I�  ���=u���?FK�  ����t�S'�q	! �  �Yхt�L8|�H�  dw�)t���v�#L�  l&��s���>��D�  �f�qs�g~��7�(�  �7�s���6�uE�  (���r�uv.�E,�  t��]r��L��v�O�  ��r��Ț�p�  �&��q�C �"5�F�  ��zIq�o����O�  �j�p�����O�  |�W�p�Ȯ�/N�  �#D5p�O���/3N�  �^�o��I��!�  `1�n��D�CE�  "Bn��u
^!E�  �WΉm����--�0�  ����l��N���pC�  P&`l����J�  �$ak�����N��  8x�j��[-=�  8R��i�y��~� �  �La8i�[�٬zF+�  �g�h�k<��@8K�  H���g�}7�ڒ�%�  ��g�mg�1&�3�   {4Wf����I�8�  �e�}�O���A�  8ӌ�d��_\���M�  P�4.d�ó�6D�  @��uc����2�I�  ��{�b��T�W�B�  `b��.�r�}�  X]�La��6MŞr<�  ��P�`���;ƥI�  p�η_��v�<�-�  �U�F^������9M�  ��\����̢N�  ��3e[��ݻ�k>?�   #J�Y�&�-D�  P�Z�X�m��4�I@�  @7eW��O���/�  �j�U���I�l�N�  �Ai0T��Wq�uI�  ��b�R��|m�:K�  �@VNQ�?|G¾d0�  `7��O�8��4�� �  �fX�L��z��B7C�  ��I�p4"%��H�  `/�G��:�
�WI�  `ȃ1D�/��!H�  @�%OA���A�9"I�  ��x�<�u*�6"dм  �7�xG��@�  @��O1���O(�;>�  ��'��8R�ؔN�   ;��*�2]��                   @G�?   �E�?   @D�?    C�?   �A�?    @�?   �>�?   @=�?   �;�?   @:�?   �8�?   �7�?    6�?   �4�?    3�?   �1�?   @0�?   �.�?   @-�?   �+�?   �*�?    )�?   �'�?    &�?   �$�?   @#�?   �!�?   @ �?   ��?   ��?    �?   ��?    �?   ��?   @�?   ��?   @�?   ��?   ��?    �?   ��?    �?   �
�?   @	�?   ��?   @�?    �?   ��?    �?   � �?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   ���?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   ���?   ���?    ��?   @��?   ��?   �~�?    ~�?   @}�?   �|�?    |�?   @{�?   �z�?   �y�?    y�?   @x�?   �w�?   �v�?   @v�?   �u�?   �t�?    t�?   @s�?   �r�?   �q�?    q�?   @p�?   �o�?    o�?   @n�?   �m�?   �l�?    l�?   @k�?   �j�?    j�?   @i�?   �h�?   �g�?    g�?   @f�?   �e�?   �d�?    d�?   �c�?   �b�?    b�?   @a�?   �`�?   �_�?    _�?   @^�?   �]�?    ]�?   @\�?   �[�?   �Z�?    Z�?   @Y�?   �X�?   �W�?    W�?   �V�?   �U�?    U�?   @T�?   �S�?   �R�?    R�?   @Q�?   �P�?    P�?   @O�?   �N�?   �M�?    M�?   @L�?   �K�?   �J�?   @J�?   �I�?   �H�?    H�?   @G�?                           �  �>Y� �"G=   � �>.ܶlW�E=   � �>jۋ�bH=     �>��^IL#=   � �>��(i�&I=   h��>g�ݟP'E=   p �>��*)��D=   � �>�&��N=   x �>.;ĝ��@=   H	 �>Qy�u�3=   �
��>�c���-=   �@�>R�ݡ�:==   ���>	��{M=    	@�>�����C=   `
��>b��ߔB=   � �>�td�C=   $��>���9��O=   � �>B� N��C=   ���>�j�&��==   ��>���.�<=    @�>`l�r�G=   ��>!���ls1=   � ?��8��=   �@?� �mN=   & ?��Ut�Q$=   X�?PiB�{^C=   ��?Gv�7��2=   �@?q�l��m+=   �?!�.j7�/=   d�?�L ��C=   �`?�m���	+=   P ?5Od%�	=   ��?�r����<   (�?*�Hga�2=   �@	?�C���I=   r 
?��s���A=   *�
?�GTi�A=   � `?�K�Ջ�D=   r" ?�Dp�`q=   L$�?��~���G=   4&�?����D=   �'@?�����E=   �) ?'P���<   �+�?f�4±cC=   �@?qW�n{;=   ��?�gC �i8=   ��?X�K�D=   P?G;��R"=   7�?�8΁3<L=   a?�rF҈K=   ^`?�_U�N=   ��?�;T��6=   � ?Ԛ����<   !�?q�W*#M=   ""�?�j�
�\M=   p#0?|I7Z#�/=   �$�?^��aDJ=   &�?��>,'1D=   B'@?�:�+NB=   �(�?�1z��@J=   * ?������3=   �+`?w�U4?�=   �,�?D��O=   ;.?$�b�� =   �/p?g)([|X>=   H1�?�>gV��=   �20?O�B��O=   *4�?bP�A��<   �5�?��e��4=   f7@?|[{�~*L=   9�?���ٹE=   t:�?G]����C=   '<P?�{m�u!K=   �=�?�
v\��4=   �??�����n=   fAp?�{7�!�O=   �B�?����=   �D ?�=u� �<=   �F�?�i&��-=   lH�?��o���N=   �I0?IT$7�QN=   �K�?Н��\�0=   �M�?0tЗ�I=   �OP?
�'��C=   uQ�?��4%@�@=   vS ?*�
qw�G=   ~U`?K ᴽ+=   �W�?F�Pn;�M=  ��, ?�]���K=  ��-8 ?�ƎI��M=  ��.h ?�5�m�3=   �/� ?�� ��M=   �0� ?�����I=   �1� ?�"���I=   �2 !?��y�$=  �4P!?�_	�D=  �.5�!?]��u�E:=  �"6�!?l�#�5=   J7�!?,����A=   u8"?��!y##�<  ��98"?�x�y�F=  ��:h"?bCڝ�D=   �;�"?u��RF=   =�"?2���w}=  �D>�"?�@(�6F=  ��? #?�'���A=   �@H#?43��A=  ��Ax#?uN}*�J=  �C�#?)�r7Yr7=  �]D�#?�.K="=   rE $?���r�=  ��F0$?3=1�Z1=   H`$?h|��=G=   gI�$?��ܩN�:=   �J�$?�4e��6=   �K�$?��{�<�9=  �=M%?uY�Pw�H=  ��NH%?��-*�8=  �Px%?�y�F�.=  �-Q�%?\9�;,=   �R�%?2�9Z�d@=   T &?~YK|=  �sU0&?WĻ��(J=  ��VX&?�R��IG=   X�&?W�	N=   �Y�&?�g�'9=   [�&?D�"^=   ���2)��$�   ����7�b�m�L�   Mӿ������(�   	ԏ��S��4�   ��_��	>��L�   |�/�����dM�   4���g±�8�   ����2�qڜ1�   �ן�qa�P�C�   Q�o�� ��%;9�   �?��_�0�C�   w��4g%6�L�   &���M��;k�@�   �ڿ�8�1�A�B�   ۏ�1�uB��   )�_����Y���   ��/�󓎣,:�   x����.Ճ^�-�   ������?�   �ޯ���ԝ�I�   -���:]=O>�   ��O�#w_jُB�   n�����(+E �   ���-�V~|_�   ����B}�_A�   C��K!ܨ�Y:�   ��_�5��G�   t�/��C���$>�   �����#���H�   m����-�
��M�   ���V���n@�   ���QU^�tA�   $�O��Ä�   ���þ��i�M�   @���K�8�|;2�   ���@�(�A�   V�����64�   ��o��ꬠTC�   9�?�&u����.�   ���~F�s:4�   �Կ��	��J�   ��_���L�II�   ����=�@�0(�   �ן��$�.�G��   ��?�}�3Rʏ3�   ����!|.4���   *ڟ�඄}��3�   �?�G"jm
>;�   ����*����O�   ���0 �:�O�   ������2K�;�   �޿�Q`���4�   ��_�� �ZD�   ���
���6�9�   *�
�����F�   �_
�T3ʢ�K�   ���	��M.�֢>�   ��	�@��_��@�   ��?	�1�\hU�   X������p�M�   &����J��x3�   ����Ҭ���   ���x�/h7�   8��L��v]E�   ����V���3�   ����B�v9�   r�_��c���M�   *����5&�L�   ���q����3�   ��?�:�R��$�   @���܎�$=�   ���K���'�   \�?��Ъ{�b>�   �����$E�vC�   ���I�w8�R'�   F��G�_j�,)�   ����+j�B�D�   |�_�`k�A�   ���%'r�BL�   ���	�T��E�   �_���GO�   ��� ��#i��#�    �� �;��^طH�   ��? �6(`J��J�   \����HB�5�   `����`��.11�   \�?��Q���D�   T����<VD��=�   D���Mϲk:UG�   ��?���,'��   �����h���UF�   ����U���ȘI�   �����t��@�5�   X�?��󕕠�4�   $������c��G�   ����y��/�C�   ������t�TM�   h�?���A�)E�   �����z�cϨN�   �����{���-��   <�?��G�#�?F�   ���}-w��F�   ����w���j'�   ���Q�x��   ��?����*
<�   4����	�,�   p��~ܾUY =�   �����˚�G�   ��쾂���p�7�   ���m�8�1<�   ����'����mN�   ��辙����L�   h���K��Y0�2�    ��̟q����   ���㾭v�Bfe9�   0���%��2�F�   ���ΥE��8�   ���߾�`�=�?�   ���ܾ��E=|
�   ���پu�M���   @��־��9��>�   ���Ӿ���9�6�   ���оk<
�xE�    ��˾�CqTR;�   ���Ǿ����dG�    �����G��gL�   @����_h�%?�   ������SS�@�                ��b��?�Wd���y>c��*GP��AiFC.ֿ      �?        53��=�?�͸�)a�<a�w>�,�?][S��q��n�C�?n�w���t�ӰY�?e�u��s�<���)kp�?&<��ߑ��țuE��?���K��a<����>��?5a1xH�<��lX��?
a�J.��<�Gr+���?qO���<���2���?R{�':@<���f��?{�N��k�Q[��?9�D9Ŗ��1l��*�?ǥl��Q��-���B�?�6�/��Q��ȘZ�?	��j@�<{Q}<�r�?u�׹A���ꍌ8���?k��#��u�o�[��?�hI{L[�<�\���?�.5�S����h1���?<d� n�<��"P��?��{�ߑ�֌b�;�?��J�uǍ<��}�I�?��~��<8bunz8�?rǶ~��<?��O�Q�?����U��<�|�eEk�?��@�3��<�c��߄�?}?�:L��������?U����<������?�8��
A�䦅��?�A�TG�<V/>����?�#�E�q<�1
��?�1�j�<1�L�p!�?|�眊<�d�<�?�Y6�!'�<�_�V�?(FN\�\��˩:7�q�?��B��:��f�m���?��<�������4ۧ�?��a�6�u���-��?�)]7����"4L���?���	ڊ<��E��?��V�#З�*.�!
�?x�0i�^���P��1�?�y_��ǁ�-�a`N�?π�z�H<W �Aj�?v�d�K��<�<�����?�b����s<����*��?V���b˙<'*6�ڿ�?�B쯗C}<������?3xj���<�,�v���?�WY�	���BfϢ��?i�v���O�V+4�?�<��z���]ʤQ�?����h���'�6Go�?��,��<�Ǘ���?��[ᕂ<)TH���?�GFL2�<�FY�&��?��i�K<<H!�o��?]�0���<	�v���?G�V�B⓼�U:�~$�?��@~���� ��4FC�?2��u<H��%"U�8b�?3Y�	���s�L�U��?d>�D�8`<�;f���?Ud�4ݛ���u��?�gV�r�/e<���?��<h:�k���Q�}��?��%<��t_��u�?�z��Gn��t��H�?�?;�el٨���gBV�_�?�m1WY$��?]�Oi��?,
�f�<��s��?/��w��2�0���?�M�L�<bN�6���?~y�]p<>T'�?*�mb�|���L��%�?�2�L����#FG�?��A��ֈ��D��h�?��ԛ�Ɵ��f��Ǌ�?:�|��<۠*B��?&K�V��<�D�2��?���2^�p�6w����?l��̅<���[�?#%X.y֝���Ͱ77�?�~���_g�R��DZ�?9�|Kv�PNޟ�}�?Ѕ|[����p��?2�Α�s���𣂑��?��q�F||<##�c��?nL�x�$x<e�]{f�?2�]IY��3-J�0�?�6�}\0�<]%>�U�?�A��n/��X�0�y�?�c��~˛<��yUk��?1�����<z�ӿk��?�l��4�����Z����?��]4͡�<f��)�?$�L�ޛ��O��3�?ׄ0^�b�:Y�rY�?�m���q��G^��v�?:�T~OXu�J�0���?.)T������K���?��-z�=�<	�[���?r�k?�����R�ݛ�?�HP�e�<z��_�@�?
ƃ�7E�<K�W.�g�?�<H�M��<���m��?D\�H��q<i��� ��?�I���u<��]U��?r��S;؍�|�J-�?�zyC7�����/�?w��q{H������X�?7[��<�����?�������2���?2�mi #�<`��!��?��xWڒ<_�{3���?[KOͥ��)��F&�?�z�'����?��.P�?�̩����<�L��Qz�?��"Ւ<ڐ�����?�(�#����g�-H��?���󓜼'Za���?�����ǝ<��k7+%�?C�����<@En[vP�?���-�ә<����{�?	5����ؐ�����?���SH�<�q�+���?�ye�t�b<      8C      8C������ ������       �?      �?��������������1g���U?���k�?wN�o���?�ł����?�9��B.�?   �����   @G��     �      �      ��       �      ��      �             ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �?5�h!���>@�������             ��      �@      �                            (   (   t b - > t m _ w d a y   > =   0   )   & &   (   t b - > t m _ w d a y   < =   6   )   )                         (   (   t b - > t m _ m d a y   > =   1   )   & &   (   (   (   _ d a y s [   t b - > t m _ m o n   +   1   ]   -   _ d a y s [   t b - > t m _ m o n   ]   )   > =   t b - > t m _ m d a y   )   | |   (   (   I S _ L E A P _ Y E A R (   t b - > t m _ y e a r   +   1 9 0 0   )   )   & &   (   t b - > t m _ m o n   = =   1   )   & &   (   t b - > t m _ m d a y   < =   2 9   )   )   )   )                                                                                     (   (   t b - > t m _ s e c   > =   0   )   & &   (   t b - > t m _ s e c   < =   5 9   )   )                           (   (   t b - > t m _ m i n   > =   0   )   & &   (   t b - > t m _ m i n   < =   5 9   )   )                           (   (   t b - > t m _ h o u r   > =   0   )   & &   (   t b - > t m _ h o u r   < =   2 3   )   )                       (   (   t b - > t m _ m o n   > =   0   )   & &   (   t b - > t m _ m o n   < =   1 1   )   )                       (   t b - > t m _ y e a r   > =   0   )             (   t b   ! =   N U L L   )         (   s i z e I n C h a r s   > =   _ A S C B U F S I Z E   )                 a s c t i m e _ s       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ a s c t i m e . c                         (   b u f f e r   ! =   N U L L   )   & &   (   s i z e I n C h a r s   >   0   )                   f:\dd\vctools\crt_bld\self_x86\crt\src\asctime.c            _ g e t _ t i m e z o n e ( & t i m e z o n e )             _ g e t _ d s t b i a s ( & d s t b i a s )             _ g e t _ d a y l i g h t ( & d a y l i g h t )             (   p t i m e   ! =   N U L L   )           _ l o c a l t i m e 6 4 _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l o c t i m 6 4 . c                       (   p t m   ! =   N U L L   )                         8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?\3&���-DT�!	�\3&��<-DT�!	@       �           �����   �����    ���                UUUUUUſ333333���m۶mۦ�颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?      �?       �9��B.�@  ׽2b      �              �7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    runtime error       
  TLOSS error
   SING error
    DOMAIN error
      R6034
An application has made an attempt to load the C runtime library without using a manifest.
This is an unsupported way to load Visual C++ DLLs. You need to modify your application to build with a manifest.
For more information, see the "Visual C++ Libraries as Shared Side-by-Side Assemblies" topic in the product documentation.
                                                                        R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
                                                  R6032
- not enough space for locale information
              R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
                      R6030
- CRT not initialized
          R6028
- unable to initialize heap
        R6027
- not enough space for lowio initialization
            R6026
- not enough space for stdio initialization
            R6025
- pure virtual function call
           R6024
- not enough space for _onexit/atexit table
            R6019
- unable to open console device
            R6018
- unexpected heap error
        R6017
- unexpected multithread lock error
            R6016
- not enough space for thread data
             
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
                               R6009
- not enough space for environment
         R6008
- not enough space for arguments
           R6002
- floating point support not loaded
            Microsoft Visual C++ Runtime Library        s t r c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   r t e r r s [ t b l i n d x ] . r t e r r t x t )                                         s t r c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   " \ n \ n " )                             ...     s t r n c p y _ s ( p c h ,   p r o g n a m e _ s i z e   -   ( p c h   -   p r o g n a m e ) ,   " . . . " ,   3 )                             <program name unknown>          s t r c p y _ s ( p r o g n a m e ,   p r o g n a m e _ s i z e ,   " < p r o g r a m   n a m e   u n k n o w n > " )                           Runtime Error!

Program:        s t r c p y _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   " R u n t i m e   E r r o r ! \ n \ n P r o g r a m :   " )                                       _ N M S G _ W R I T E           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c r t 0 m s g . c                         s t r n c p y _ s ( * s t r a d d r e s s ,   o u t s i z e ,   p c b u f f e r ,   o u t s i z e   -   1 )                         _ _ g e t l o c a l e i n f o               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t h e l p . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\inithelp.c           f:\dd\vctools\crt_bld\self_x86\crt\src\osfinfo.c            _ g e t _ o s f h a n d l e             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o s f i n f o . c                         f:\dd\vctools\crt_bld\self_x86\crt\src\ioinit.c             _ _ l o c t o t i m e 6 4 _ t               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d t o x t m 6 4 . c                       _ o p e n       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o p e n . c                       ( p a t h   ! =   N U L L )             ( ( p m o d e   &   ( ~ ( _ S _ I R E A D   |   _ S _ I W R I T E ) ) )   = =   0 )                     _ s o p e n _ h e l p e r           ( p f h   ! =   N U L L )           0   & &   " O n l y   U T F - 1 6   l i t t l e   e n d i a n   &   U T F - 8   i s   s u p p o r t e d   f o r   r e a d s "                               0   & &   " I n t e r n a l   E r r o r "           ( o f l a g   &   ( _ O _ T E X T   |   _ O _ W T E X T   |   _ O _ U 1 6 T E X T   |   _ O _ U 8 T E X T )   )   ! =   0                           (   " I n v a l i d   s h a r i n g   f l a g "   ,   0   )                 (   " I n v a l i d   o p e n   f l a g "   ,   0   )               _ g e t _ f m o d e ( & f m o d e )             _ t s o p e n _ n o l o c k         _ w o p e n     _ w s o p e n _ h e l p e r                   �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��                    tan cos sin modf    floor   ceil    atan    exp10   acos    asin    pow exp log10   log                                           �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      �                                                                                                                                                                                                                                                                                                                                                                                                                                                            s t r c p y _ s ( * e n v ,   c c h a r s ,   p )               _ s e t e n v p             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t d e n v p . c                         f:\dd\vctools\crt_bld\self_x86\crt\src\stdenvp.c            f:\dd\vctools\crt_bld\self_x86\crt\src\stdargv.c            f:\dd\vctools\crt_bld\self_x86\crt\src\a_env.c          f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ h e a p i n i t . c                       _ c r t h e a p           �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �                               ( " i n c o n s i s t e n t   I O B   f i e l d s " ,   s t r e a m - > _ p t r   -   s t r e a m - > _ b a s e   > =   0 )                             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f l s b u f . c                         s t r   ! =   N U L L       ( n u l l )     (null)             EEE50 P    ( 8PX 700WP        `h````  xpxxxx                          f:\dd\vctools\crt_bld\self_x86\crt\src\output.c             ( " ' n '   f o r m a t   s p e c i f i e r   d i s a b l e d " ,   0 )                 ( c h   ! =   _ T ( ' \ 0 ' ) )         _ o u t p u t _ l       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o u t p u t . c                           ( " M i s s i n g   p o s i t i o n   i n   t h e   f o r m a t   s t r i n g " ,   0 )                         ( ( s t a t e   = =   S T _ N O R M A L )   | |   ( s t a t e   = =   S T _ T Y P E ) )                         _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ l o n g _ l o n g _ a r g ,   c h ,   f l a g s )                                 _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ i n t 6 4 _ a r g ,   c h ,   f l a g s )                                 p a s s   = =   F O R M A T _ O U T P U T _ P A S S             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ d o u b l e _ a r g ,   c h ,   f l a g s )                               _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ p t r _ a r g ,   c h ,   f l a g s )                             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ s h o r t _ a r g ,   c h ,   f l a g s )                                 ( ( t y p e _ p o s > = 0 )   & &   ( t y p e _ p o s < _ A R G M A X ) )                       _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ p r e c i s _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                                 ( ( p r e c i s _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                     _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ w i d t h _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                                   ( ( w i d t h _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                       ( " I n c o r r e c t   f o r m a t   s p e c i f i e r " ,   0 )                       ( ( t y p e _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                 _ o u t p u t _ p _ l           �������             ��      �@      �                    f:\dd\vctools\crt_bld\self_x86\crt\src\_sftbuf.c            f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ s f t b u f . c                         f l a g   = =   0   | |   f l a g   = =   1             f w r i t e     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f w r i t e . c                           ( " I n c o n s i s t e n t   S t r e a m   C o u n t .   F l u s h   b e t w e e n   c o n s e c u t i v e   r e a d   a n d   w r i t e " ,   s t r e a m - > _ c n t   > =   0 )                                         n u m   < =   ( S I Z E _ M A X   /   s i z e )             ( b u f f e r   ! =   N U L L )         _ f w r i t e _ n o l o c k         _ f i l e n o       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f i l e n o . c                       ( _ o s f i l e ( f i l e d e s )   &   F O P E N )             _ c o m m i t       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c o m m i t . c                           ( f i l e d e s   > =   0   & &   ( u n s i g n e d ) f i l e d e s   <   ( u n s i g n e d ) _ n h a n d l e )                         _ w r i t e     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w r i t e . c                     i s l e a d b y t e ( _ d b c s B u f f e r ( f h ) )               ( ( c n t   &   1 )   = =   0 )         _ w r i t e _ n o l o c k           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ h a n d l e r . c p p                         p n h   = =   0         Assertion Failed    Error   Warning     `VXVDV    _ C r t S e t R e p o r t H o o k 2             Microsoft Visual C++ Debug Library          Debug %s!

Program: %s%s%s%s%s%s%s%s%s%s%s%s

(Press Retry to debug the application)                    
Module:    
File:      
Line:      Expression:         

For information on how your program can cause an assertion
failure, see the Visual C++ documentation on asserts.                              s t r c p y _ s ( s z E x e N a m e ,   2 6 0 ,   " < p r o g r a m   n a m e   u n k n o w n > " )                         _ _ c r t M e s s a g e W i n d o w A           _ e x p a n d _ b a s e             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ e x p a n d . c                       p B l o c k   ! =   N U L L         HeapQueryInformation        k e r n e l 3 2 . d l l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s b h e a p . c                           ( t h r e s h o l d   < =   M A X _ A L L O C _ D A T A _ S I Z E )   & &   _ _ s b h _ h e a p _ i n i t ( t h r e s h o l d )                             _ s e t _ s b h _ t h r e s h o l d                 t h r e s h o l d   < =   M A X _ A L L O C _ D A T A _ S I Z E                 _ s e t _ a m b l k s i z           0   <   s i z e   & &   s i z e   < =   U I N T _ M A X                 _ g e t _ a m b l k s i z           p S i z e   ! =   N U L L           f:\dd\vctools\crt_bld\self_x86\crt\src\mbctype.c            LC_TIME     LC_NUMERIC      LC_MONETARY     LC_CTYPE    LC_COLLATE      LC_ALL  �\    ߯p\�V��d\�V�T\�VБD\�Vf�8\�V��                	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~                         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s e t l o c a l . c                       ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w l o c a l e   ! =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w r e f c o u n t   ! =   N U L L ) )   | |   ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w l o c a l e   = =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w r e f c o u n t   = =   N U L L ) )                                                                                         _ c o n f i g t h r e a d l o c a l e           ( " I n v a l i d   p a r a m e t e r   f o r   _ c o n f i g t h r e a d l o c a l e " , 0 )                       f:\dd\vctools\crt_bld\self_x86\crt\src\setlocal.c           s e t l o c a l e       L C _ M I N   < =   _ c a t e g o r y   & &   _ c a t e g o r y   < =   L C _ M A X                     s t r n c p y _ s ( l c t e m p ,   ( s i z e o f ( l c t e m p )   /   s i z e o f ( l c t e m p [ 0 ] ) ) ,   s ,   l e n )                               _ s e t l o c a l e _ n o l o c k           ;   =;  s t r c p y _ s ( p c h   +   s i z e o f ( i n t ) ,   c c h   -   s i z e o f ( i n t ) ,   l c t e m p )                         _ s e t l o c a l e _ s e t _ c a t             s t r c a t _ s ( p c h ,   c c h ,   " ; " )               _ s e t l o c a l e _ g e t _ a l l             =       s t r c p y _ s ( o u t p u t ,   s i z e I n C h a r s ,   c a c h e o u t )                   s t r n c p y _ s ( c a c h e i n ,   c a c h e i n S i z e ,   s o u r c e ,   c h a r a c t e r s I n S o u r c e   +   1 )                               C   s t r c p y _ s ( o u t p u t ,   s i z e I n C h a r s ,   " C " )                 _ e x p a n d l o c a l e           s t r c a t _ s ( o u t s t r ,   s i z e I n B y t e s ,   (   * ( c h a r   *   * ) ( ( s u b s t r   + =   (   ( s i z e o f ( c h a r   * )   +   s i z e o f ( i n t )   -   1 )   &   ~ ( s i z e o f ( i n t )   -   1 )   ) )   -   (   ( s i z e o f ( c h a r   * )   +   s i z e o f ( i n t )   -   1 )   &   ~ ( s i z e o f ( i n t )   -   1 )   ) )   ) )                                                                           _ s t r c a t s             s t r n c p y _ s ( n a m e s - > s z C o d e P a g e ,   ( s i z e o f ( n a m e s - > s z C o d e P a g e )   /   s i z e o f ( n a m e s - > s z C o d e P a g e [ 0 ] ) ) ,   l o c a l e ,   l e n )                                               s t r n c p y _ s ( n a m e s - > s z C o u n t r y ,   ( s i z e o f ( n a m e s - > s z C o u n t r y )   /   s i z e o f ( n a m e s - > s z C o u n t r y [ 0 ] ) ) ,   l o c a l e ,   l e n )                                             s t r n c p y _ s ( n a m e s - > s z L a n g u a g e ,   ( s i z e o f ( n a m e s - > s z L a n g u a g e )   /   s i z e o f ( n a m e s - > s z L a n g u a g e [ 0 ] ) ) ,   l o c a l e ,   l e n )                                           _., s t r n c p y _ s ( n a m e s - > s z C o d e P a g e ,   ( s i z e o f ( n a m e s - > s z C o d e P a g e )   /   s i z e o f ( n a m e s - > s z C o d e P a g e [ 0 ] ) ) ,   & l o c a l e [ 1 ] ,   1 6 - 1 )                                             _ _ l c _ s t r t o l c         .   _   s t r c p y _ s ( l o c a l e ,   s i z e I n B y t e s ,   ( c h a r   * ) n a m e s - > s z L a n g u a g e )                         _ _ l c _ l c t o s t r         s p r i n t f           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s p r i n t f . c                         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i s c t y p e . c                         ( u n s i g n e d ) ( c   +   1 )   < =   2 5 6             MSPDB80.DLL     r   PDBOpenValidate5    EnvironmentDirectory        SOFTWARE\Microsoft\VisualStudio\9.0\Setup\VS            RegCloseKey     RegQueryValueExA    RegOpenKeyExA   ADVAPI32.DLL    _ c o n t r o l f p _ s             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ t r a n \ c o n t r l f p . c                           ( " I n v a l i d   i n p u t   v a l u e " ,   0 )             p f l t   ! =   N U L L         s i z e I n B y t e s   >   ( s i z e _ t ) ( ( d i g i t s   >   0   ?   d i g i t s   :   0 )   +   1 )                           _ f p t o s t r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f p t o s t r . c                       s t r c p y _ s ( r e s u l t s t r ,   r e s u l t s i z e ,   a u t o f o s . m a n )                     _ f l t o u t 2             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ c f o u t . c                         _ s e t _ o u t p u t _ f o r m a t             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o u t p u t f o r m a t . c                               ( o p t i o n s   &   ~ _ T W O _ D I G I T _ E X P O N E N T )   = =   0                    Complete Object Locator'        Class Hierarchy Descriptor'         Base Class Array'       Base Class Descriptor at (          Type Descriptor'       `local static thread guard'         `managed vector copy constructor iterator'          `vector vbase copy constructor iterator'            `vector copy constructor iterator'          `dynamic atexit destructor for '        `dynamic initializer for '      `eh vector vbase copy constructor iterator'         `eh vector copy constructor iterator'           `managed vector destructor iterator'        `managed vector constructor iterator'           `placement delete[] closure'        `placement delete closure'      `omni callsig'       delete[]    new[]  `local vftable constructor closure'         `local vftable'     `RTTI   `EH `udt returning'     `copy constructor closure'      `eh vector vbase constructor iterator'          `eh vector destructor iterator'         `eh vector constructor iterator'        `virtual displacement map'      `vector vbase constructor iterator'         `vector destructor iterator'        `vector constructor iterator'       `scalar deleting destructor'        `default constructor closure'       `vector deleting destructor'        `vbase destructor'      `string'    `local static guard'        `typeof'    `vcall'     `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ()  >=  >   <=  <   %   ->* &   +   --  ++  *   ->  operator    []  !=  ==  !   <<  >>   delete      new    __unaligned     __restrict      __ptr64     __clrcall   __fastcall      __thiscall      __stdcall   __pascal    __cdecl     __based(        �w�w�w�w�w�w�w�wtwdwLr�q�q�q�q\wPw8cLwHwDw@w<w8w,w(w$w ww�-www0www w�v\N�v`V�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�vtvhvPv,vv�u�u�upuPu(u u�t�t�t�t�t|tPtHt<t(tt�s�s�sXs$ss�r�r|rHr$rL                                                                            CV:     ::  '   `   generic-type-   template-parameter-     ''  `anonymous namespace'       `non-type-template-parameter        `template-parameter     void    NULL    extern "C"      [thunk]:    public:     protected:      private:    virtual     static      `template static data member destructor helper'             `template static data member constructor helper'            `local static destructor helper'        `adjustor{      `vtordisp{      `vtordispex{    }'  }'  )   void    volatile    ,<ellipsis>     ,...    <ellipsis>       throw(      volatile   const   signed      unsigned    UNKNOWN     __w64   wchar_t     __int128    __int64     __int32     __int16     __int8  bool    double  long    float   long    int short   char    enum    cointerface     coclass     class   struct      union   `unknown ecsu'      int     short   char    const   volatile    cli::pin_ptr<   cli::array<     )[  {flat}  s   {for    ,�,�,�    f��י    ����    '���a�    ���݉     ??     ����    _ m b s t o w c s _ l _ h e l p e r                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b s t o w c s . c                       s   ! =   N U L L       r e t s i z e   < =   s i z e I n W o r d s             b u f f e r S i z e   < =   I N T _ M A X           _ m b s t o w c s _ s _ l           ( p w c s   = =   N U L L   & &   s i z e I n W o r d s   = =   0 )   | |   ( p w c s   ! =   N U L L   & &   s i z e I n W o r d s   >   0 )                                   ( L " S t r i n g   i s   n o t   n u l l   t e r m i n a t e d "   & &   0 )                   S t r i n g   i s   n o t   n u l l   t e r m i n a t e d               s t r c a t _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s c a t _ s . i n l                           ( c o u n t   = =   0 )   | |   ( s t r i n g   ! =   N U L L )                 _ v s n p r i n t f _ h e l p e r           ( " B u f f e r   t o o   s m a l l " ,   0 )               s t r i n g   ! =   N U L L   & &   s i z e I n B y t e s   >   0                   _ v s p r i n t f _ s _ l           f o r m a t   ! =   N U L L         _ v s n p r i n t f _ s _ l         l e n g t h   <   s i z e I n T C h a r s           2   < =   r a d i x   & &   r a d i x   < =   3 6                   s i z e I n T C h a r s   >   ( s i z e _ t ) ( i s _ n e g   ?   2   :   1 )                   s i z e I n T C h a r s   >   0         x t o a _ s     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ x t o a . c                       x 6 4 t o a _ s         _ w c s t o m b s _ l _ h e l p e r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c s t o m b s . c                       p w c s   ! =   N U L L         s i z e I n B y t e s   >   r e t s i z e           _ w c s t o m b s _ s _ l           ( d s t   ! =   N U L L   & &   s i z e I n B y t e s   >   0 )   | |   ( d s t   = =   N U L L   & &   s i z e I n B y t e s   = =   0 )                               w c s c a t _ s         _ v s w p r i n t f _ h e l p e r               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v s w p r i n t . c                       s t r i n g   ! =   N U L L   & &   s i z e I n W o r d s   >   0                   _ v s w p r i n t f _ s _ l         _ v s n w p r i n t f _ s _ l           x t o w _ s     x 6 4 t o w _ s         SystemFunction036       ( " r a n d _ s   i s   n o t   a v a i l a b l e   o n   t h i s   p l a t f o r m " ,   0 )                       r a n d _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ r a n d _ s . c                       _ R a n d o m V a l u e   ! =   N U L L             _ w o u t p u t _ l         _ v s w p r i n t f _ l         _ v s c w p r i n t f _ h e l p e r             SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec                _ g e t _ d a y l i g h t               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t i m e s e t . c                         ( _ D a y l i g h t   ! =   N U L L )           _ g e t _ d s t b i a s         ( _ D a y l i g h t _ s a v i n g s _ b i a s   ! =   N U L L )                 _ g e t _ t i m e z o n e           ( _ T i m e z o n e   ! =   N U L L )           _ I n d e x   = =   0   | |   _ I n d e x   = =   1             _ R e t u r n V a l u e   ! =   N U L L             _ g e t _ t z n a m e           ( _ B u f f e r   ! =   N U L L   & &   _ S i z e I n B y t e s   >   0 )   | |   ( _ B u f f e r   = =   N U L L   & &   _ S i z e I n B y t e s   = =   0 )                                   s t r n c p y _ s ( t z n a m e [ 1 ] ,   6 4 ,   T Z ,   3 )                   s t r n c p y _ s ( t z n a m e [ 0 ] ,   6 4 ,   T Z ,   3 )                   s t r c p y _ s ( l a s t T Z ,   s t r l e n ( T Z )   +   1 ,   T Z )                 f:\dd\vctools\crt_bld\self_x86\crt\src\tzset.c          TZ  _ t z s e t _ n o l o c k           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t z s e t . c                     _ i s i n d s t _ n o l o c k           c v t d a t e       _ g m t i m e 6 4 _ s       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ g m t i m e 6 4 . c                       _ g m t i m e 3 2 _ s           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ g m t i m e . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\gmtime.c             _ s e t _ e r r o r _ m o d e           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ e r r m o d e . c                         ( " I n v a l i d   e r r o r _ m o d e " ,   0 )               GetUserObjectInformationA       MessageBoxA     USER32.DLL      s t r n c p y _ s       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s n c p y _ s . i n l                         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m a l l o c . h                           ( " C o r r u p t e d   p o i n t e r   p a s s e d   t o   _ f r e e a " ,   0 )                   _ l s e e k i 6 4           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l s e e k i 6 4 . c                       ( s i z e   > =   0 )       _ c h s i z e _ s           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c h s i z e . c                       ( c n t   < =   I N T _ M A X )         _ r e a d           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ r e a d . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\read.c           ( i n p u t b u f   ! =   N U L L )             _ r e a d _ n o l o c k         _ l s e e k     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l s e e k . c                     ( " I n v a l i d   f i l e   d e s c r i p t o r " , 0 )               _ s e t m o d e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s e t m o d e . c                         ( ( m o d e   = =   _ O _ T E X T )   | |   ( m o d e   = =   _ O _ B I N A R Y )   | |   ( m o d e   = =   _ O _ W T E X T )   | |   ( m o d e   = =   _ O _ U 8 T E X T )   | |   ( m o d e   = =   _ O _ U 1 6 T E X T ) )                                               _ s e t _ f m o d e         ( ( m o d e   = =   _ O _ T E X T )   | |   ( m o d e   = =   _ O _ B I N A R Y )   | |   ( m o d e   = =   _ O _ W T E X T ) )                             _ g e t _ f m o d e         ( p M o d e   ! =   N U L L )           _nextafter      _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh    f:\dd\vctools\crt_bld\self_x86\crt\src\_getbuf.c            f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ g e t b u f . c                         _ i s a t t y           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i s a t t y . c                       p r i n t f         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ p r i n t f . c                       _ w c t o m b _ s _ l       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c t o m b . c                       s i z e I n B y t e s   < =   I N T _ M A X                 i b a s e   = =   0   | |   ( 2   < =   i b a s e   & &   i b a s e   < =   3 6 )                   s t r t o x l       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r t o l . c                       n p t r   ! =   N U L L             ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp                       _ o u t p u t _ s _ l       f c l o s e     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f c l o s e . c                       _ f c l o s e _ n o l o c k         ( s t r   ! =   N U L L )           _ c p u t w s       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ p u t w c h . c                           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b t o w c . c                           _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   1   | |   _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   2                                                                                                                                                                                                                                                                                                                                   ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t t i m e . c                       p l o c i - > l c _ t i m e _ c u r r - > r e f c o u n t   >   0                   f:\dd\vctools\crt_bld\self_x86\crt\src\inittime.c           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t n u m . c                         p l o c i - > l c o n v _ n u m _ r e f c o u n t   >   0               f:\dd\vctools\crt_bld\self_x86\crt\src\initnum.c                f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t m o n . c                         p l o c i - > l c o n v _ m o n _ r e f c o u n t   >   0               f:\dd\vctools\crt_bld\self_x86\crt\src\initmon.c            p l o c i - > c t y p e 1 _ r e f c o u n t   >   0                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t c t y p . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\initctyp.c           HH:mm:ss    dddd, MMMM dd, yyyy     MM/dd/yy    PM  AM  December    November    October     September   August  July    June    April   March   February    January     Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday     Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > w d a y [ n ] )                       s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > w d a y _ a b b r [ n ] )                         _ G e t d a y s _ l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r f t i m e . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\strftime.c               s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > m o n t h [ n ] )                     s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > m o n t h _ a b b r [ n ] )                       _ G e t m o n t h s _ l             s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > w w _ t i m e f m t )                     s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > w w _ l d a t e f m t )                           s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > w w _ s d a t e f m t )                           s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > a m p m [ 1 ] )                   s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > a m p m [ 0 ] )                   s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > m o n t h [ n ] )                         s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > m o n t h _ a b b r [ n ] )                       s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > w d a y [ n ] )                   s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > w d a y _ a b b r [ n ] )                     _ G e t t n a m e s _ l         F A L S E           ( " I n v a l i d   M B C S   c h a r a c t e r   s e q u e n c e   p a s s e d   t o   s t r f t i m e " , 0 )                         t i m e p t r   ! =   N U L L           (   f o r m a t   ! =   N U L L   )             (   m a x s i z e   ! =   0   )         _ S t r f t i m e _ l       (   s t r i n g   ! =   N U L L   )                 (   " I n v a l i d   f o r m a t   d i r e c t i v e "   ,   0   )                     (   t i m e p t r - > t m _ y e a r   > =   - 1 9 0 0   )   & &   (   t i m e p t r - > t m _ y e a r   < =   8 0 9 9   )                           (   t i m e p t r - > t m _ y e a r   > = 0   )             (   (   t i m e p t r - > t m _ s e c   > = 0   )   & &   (   t i m e p t r - > t m _ s e c   < =   5 9   )   )                         (   (   t i m e p t r - > t m _ m i n   > = 0   )   & &   (   t i m e p t r - > t m _ m i n   < =   5 9   )   )                         (   (   t i m e p t r - > t m _ y d a y   > = 0   )   & &   (   t i m e p t r - > t m _ y d a y   < =   3 6 5   )   )                           (   (   t i m e p t r - > t m _ h o u r   > = 0   )   & &   (   t i m e p t r - > t m _ h o u r   < =   2 3   )   )                             (   (   t i m e p t r - > t m _ m d a y   > = 1   )   & &   (   t i m e p t r - > t m _ m d a y   < =   3 1   )   )                             (   (   t i m e p t r - > t m _ m o n   > = 0   )   & &   (   t i m e p t r - > t m _ m o n   < =   1 1   )   )                         _ e x p a n d t i m e           (   (   t i m e p t r - > t m _ w d a y   > = 0   )   & &   (   t i m e p t r - > t m _ w d a y   < =   6   )   )                               ( " I n v a l i d   M B C S   c h a r a c t e r   s e q u e n c e   p a s s e d   i n t o   s t r f t i m e " , 0 )                             ( " I n v a l i d   M B C S   c h a r a c t e r   s e q u e n c e   f o u n d   i n   l o c a l e   A M P M   s t r i n g " , 0 )                               a/p am/pm   united-states   united-kingdom      trinidad & tobago       south-korea     south-africa    south korea     south africa    slovak  puerto-rico     pr-china    pr china    nz  new-zealand     hong-kong   holland     great britain   england     czech   china   britain     america     usa us  uk  swiss   swedish-finland     spanish-venezuela       spanish-uruguay     spanish-puerto rico     spanish-peru    spanish-paraguay    spanish-panama      spanish-nicaragua       spanish-modern      spanish-mexican     spanish-honduras    spanish-guatemala       spanish-el salvador     spanish-ecuador     spanish-dominican republic      spanish-costa rica      spanish-colombia    spanish-chile   spanish-bolivia     spanish-argentina       portuguese-brazilian        norwegian-nynorsk       norwegian-bokmal    norwegian   italian-swiss   irish-english   german-swiss    german-luxembourg       german-lichtenstein     german-austrian     french-swiss    french-luxembourg       french-canadian     french-belgian      english-usa     english-us      english-uk      english-trinidad y tobago       english-south africa        english-nz      english-jamaica     english-ire     english-caribbean       english-can     english-belize      english-aus     english-american    dutch-belgian   chinese-traditional     chinese-singapore       chinese-simplified      chinese-hongkong    chinese     chi chh canadian    belgian     australian      american-english    american english    american    ��ENU ��ENU |�ENU l�ENA `�NLB T�ENC P�ZHH L�ZHI @�CHS ,�ZHH �CHS ��ZHI ��CHT ��NLB ��ENU ��ENA ��ENL ��ENC t�ENB d�ENI P�ENJ @�ENZ $�ENS �ENT ��ENG ��ENU ��ENU ��FRB ��FRC ��FRL ��FRS p�DEA X�DEC @�DEL 0�DES  �ENI �ITS �NOR �NOR ؿNON ��PTB ��ESS ��ESB ��ESL l�ESO T�ESC 4�ESD  �ESF �ESE �ESG ܾESH ȾESM ��ESN ��ESI ��ESA t�ESZ d�ESR L�ESU 8�ESY  �ESV �SVF �DES  �ENG ��ENU ��ENU                                                                                                         �USA �GBR ؽCHN нCZE ĽGBR ��GBR ��NLD ��HKG ��NZL ��NZL |�CHN p�CHN `�PRI X�SVK H�ZAF 8�KOR (�ZAF �KOR  �TTO  �GBR �GBR ܼUSA ��USA                                     6-    Norwegian-Nynorsk           s t r c p y _ s ( l p O u t S t r - > s z L a n g u a g e ,   ( s i z e o f ( l p O u t S t r - > s z L a n g u a g e )   /   s i z e o f ( l p O u t S t r - > s z L a n g u a g e [ 0 ] ) ) ,   " N o r w e g i a n - N y n o r s k " )                                                   _ _ g e t _ q u a l i f i e d _ l o c a l e                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ g e t q l o c . c                         OCP 0   ACP  _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   n e w c t r l ,   m a s k   &   ~ 0 x 0 0 0 8 0 0 0 0 )                         _ s e t _ c o n t r o l f p         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ t r a n \ i 3 8 6 \ i e e e 8 7 . c                             _ _ s t r g t o l d 1 2 _ l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ i n c l u d e \ s t r g t o l d 1 2 . i n l                             _ L o c a l e   ! =   N U L L           1#QNAN  s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # Q N A N " )                 1#INF       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N F " )                   1#IND       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N D " )                   1#SNAN      s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # S N A N " )                 $ I 1 0 _ O U T P U T       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ x 1 0 f o u t . c                             _ w o u t p u t _ s _ l         _ w o u t p u t _ p _ l         f p u t w c     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f p u t w c . c                           ( _ t c s n l e n ( o p t i o n ,   _ M A X _ E N V )   <   _ M A X _ E N V )                   g e t e n v     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ g e t e n v . c                       ( o p t i o n   ! =   N U L L )             _ t c s n l e n ( * s e a r c h   +   l e n g t h   +   1 ,   _ M A X _ E N V )   <   _ M A X _ E N V                           s t r c p y _ s ( b u f f e r ,   s i z e I n T C h a r s ,   s t r )                   ( b u f f e r   ! =   N U L L   & &   s i z e I n T C h a r s   >   0 )   | |   ( b u f f e r   = =   N U L L   & &   s i z e I n T C h a r s   = =   0 )                                   _ g e t e n v _ s _ h e l p e r         p R e t u r n V a l u e   ! =   N U L L             s t r c p y _ s ( * p B u f f e r ,   s i z e ,   s t r )               v a r n a m e   ! =   N U L L           _ d u p e n v _ s _ h e l p e r         p B u f f e r   ! =   N U L L           v p r i n t f _ h e l p e r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v p r i n t f . c                         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f r e e b u f . c                       s t r e a m   ! =   N U L L         CONIN$  CONOUT$     f:\dd\vctools\crt_bld\self_x86\crt\src\convrtcp.c           _ s t r i c m p _ l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r i c m p . c                         _ s t r i c m p         c o u n t   < =   I N T _ M A X         _ s t r n i c m p _ l           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r n i c m p . c                       _ s t r n i c m p       s t r t o x q           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r t o q . c                       w c s t o x l       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c s t o l . c                       n   < =   I N T _ M A X         s 2   ! =   N U L L         _ m b s n b i c o l l _ l               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b s n b i c o . c                       s 1   ! =   N U L L         f:\dd\vctools\crt_bld\self_x86\crt\src\wtombenv.c           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ a _ c m p . c                     c c h C o u n t 1 = = 0   & &   c c h C o u n t 2 = = 1   | |   c c h C o u n t 1 = = 1   & &   c c h C o u n t 2 = = 0                             _ s t r i n g 2   ! =   N U L L         _ s t r n i c o l l _ l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r n i c o l . c                       _ s t r i n g 1   ! =   N U L L         s t r c p y _ s ( n a m e ,   s t r l e n ( o p t i o n )   +   2 ,   o p t i o n )                     ( " C R T   L o g i c   e r r o r   d u r i n g   s e t e n v " , 0 )                   f:\dd\vctools\crt_bld\self_x86\crt\src\setenv.c                 _ t c s n l e n ( e q u a l   +   1 ,   _ M A X _ E N V )   <   _ M A X _ E N V                     e q u a l   -   o p t i o n   <   _ M A X _ E N V               _ _ c r t s e t e n v       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s e t e n v . c                       p o p t i o n   ! =   N U L L               s t r c p y _ s ( * n e w e n v p t r ,   e n v p t r S i z e ,   * o l d e n v p t r )                     c o p y _ e n v i r o n         _ m b s c h r _ l           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b s c h r . c                       s t r i n g   ! =   N U L L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     RSDSF6Y;+�E�X��u��  C:\Program Files (x86)\CINEMA 4D R10\plugins\VRMLExporter\obj\vrmlexporter_Win32_Debug.pdb                                                                                                                                                                                                                                                                                                      @�               ,�    @�d�����    @       ����    @   �        $@       ����    @   ��                   ��    d�����    D@       ����    @   ��                   ��    ����    `@        ����    @   �                   (�    ��                $@��                D@��                �@x�               ��    ����    �@       ����    @   x�        �@        ����    @   ��                   ��    ��                �@�               (�    8�\���    �@       ����    @   �        �@       ����    @   ��                   ��    \���                �@��                A��               ��    ��d�����    A       ����    @   ��                    HA4�               H�    X�|���    HA       ����    @   4�        hA       ����    @   ��                   ��    |���    �A        ����    @   ��                   ��    ��                �A�               ,�    @�d�����    �A       ����    @   �        �A       ����    @   ��                   ��    d�����                �A��                �A��               ��     �|���    �A       ����    @   ��                    lB<�               P�    \���    lB       ����    @   <�        �B        ����    @   ��                   ��    ��                �B��                �B��               �    �    �B        ����    @   ��                    `@�                �A��                hA��                �B��               ��    ��    �B        ����    @   ��                    C��               ��    ���    C       ����    @   ��                    4CD�               X�    h����    4C       ����    @   D�                    dC��               ��    ����    dC       ����    @   ��                    �C �               �     ���    �C       ����    @    �                    D\�               p�    ��\���    D       ����    @   \�                    ,D��               ��    ��\���    ,D       ����    @   ��                    pD�               0�    8�    pD        ����    @   �                    �@��                �D��               ��    ����    �D       ����    @   ��                    �D��               ��    ���    �D       ����    @   ��                    �DD�               X�    h����    �D       ����    @   D�                    �H��               ��    ����    �H       ����    @   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍٍ                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ������    ��    á"�   ��                               ����������"�   ��                               ����`�"�   0�                           ������"�   `�                           ������"�   ��                           "�   ��                       ��������������������(�����3�����A�����L�            "�   L�                       ������������   ������������̣   ԣ   ߣ   �   ��    �   �   �   !�   ,�   7�   B�   M�   X�   c�   n�                    �����"�    �                           ����0�����;�"�   0�                               ������    ��   ��"�   l�                               ����Х    إ   �"�   ��                               ���� �"�   ��                           "�   H�                       ����`�    h�   s�   ~�    ��   ��        �����    �"�   ��                               ����@�    H�"�   ��                               ������    ��   ��"�   ��                                   �    P�       `���        �@    ����       �        �@    ����       Z�    �����"�   ��                           �����"�   ��                           ����H�    @�"�    �                               ������    ��   ��"�   <�                               �����    �"�   ��                               ����p�"�   ��                           @           �a����    ����                  ��"�   ��   �                       ����ة    Щ"�   L�                               @           �q����    ����                  ��"�   ��   ��                           
�    ,�    ����`�"�   ��                              @�`���        �@    ����    ,   $�        �@    ����    ,   L�    ������"�   ��                           ����Ъ"�   ��                           ���� �"�   ��                           ����0�"�   �                           ����`�"�   @�                           ������"�   p�                           @           ��@           (�����    ����                  "�   ��                               ��              ��                �����������"�   <                                "�#   �                        ����@�    H�    S�    ^�   f�   q�   |�   ��   ��   ��	   ��
   ��   ��   ɬ   Ԭ   ߬   �   ��    �   �   �   !�   ,�   7�   B�   M�   X�   c�   n�   y�   ��   ��   ��    ��!   ��                                ����P�    X�"�   �                               ������    ��   ��"�                                  "�   x                       ���� �    �   �   !�   ,�����7�   B�   M�   X�����c�����n�            "�                           ����Я    د   �   �   ��   �   �   �   %�   0�   ;�   F�   T�   _�                "�,   �                       ����а    ۰   �   �������   �   �   �   (�   3�	   >�
   I�   T�   _�   j�   u�������   ��   ��   ��   ��   ��   ±   ͱ   ر   �   �   �������   �   �   %�   0�    ;�!   F�"   Q�#   \�$   g�%   r�&   }�'   ��(   ��)   ��*   ��                                        ����`�    h�   s�"�   ,                               "�   �                       ������    ȳ   г   ۳   �   �   ��   �   �   �   (�
   3�   >�   I�
   T�
   _�   j�   u�   ��   ��   ��   ��   ��   ��   ´                        "�   �                       ����P�    X�   `�   h�   p�   x�   ��   ��   ��   ��	   ��
   ��   µ   ͵   ص   �   �   �   ��                    ����p�"�   D                           ������"�   t                           ����ض    ж"�   �                               ����8�    0�   W�"�   �                               ������"�   $                           "�   x                       ����з    ط   �   �   ��   
�        ����P�    X�   c�   q�"�   �                               ������"�   �                           �����    �   �   ��"�   ,	                               ����@�    K�"�   x	                               ������"�   �	                           ������    ȹ"�   �	                               ���� �    �   �"�    
                               ������    P�   X�   c�"�   d
                               �����"�   �
                           "�	                          ����F�     �   (�   0�   ;�   e�   p�   {�   ��            �����"�   X                           �����"�   �                           ����@�    H�   S�    ^�"�   �                               ������"�                              ����ؼ    м"�   4                               ����C�    0�   8�"�   p                               "�   �                       ������    ��   ��   ��   ý   ν        �����"�                              ����H�    @�"�   @                               ������"�   |                           "�   �                       ����о    ؾ   �   �   �   ��   �   �            @           �L����    ����                  "�   ,   <                       "�   �                       ������    ��   ��   ��   ��    ��        ���� �"�   �                           ����8�    0�"�                                  "�   h                       ������    ��   ��   ��   ��   �        @           �a����    ����                  �"�   �   �                       ������"�                               ������"�   0                           "�   �                       ���� �     �   �   �   �        ������"�   �                           ������    ��"�   �                               @           qp@           �n"�   �   d                           0             ���� �                    (�                  0�                ����p�"�   �                           "�   (                       ������    ��   ��   ��   ��        ���� �"�   X                           @           Љ            �"�   �   �               ����@�    H�   P�   X�   c�                 k�                @           ������    ����                   "�   0   @                       ������    ��   ��"�   �                               ����0�"�   �                           ����p�"�   �                           @           X�����    ����                  $"�   4   D                       "�   �                       ������������   ��   ��   ��        ����@�"�   �                           "�
   ,                       ����p�    x�   ��   ��   ��   ��   ��   ��   ��   ��            "�   �                       ����0�    8�   C�   N�    Y�   d�    o�    z�    ��    ��	   ��
   ��   ��   ��   ��   ��   ��   ��   ��    ��   	�   �    �   *�   5�   @�   K�   V�                            "�   �                       ������    ��   ��   ��    	�   �    �   *�   5�   @�	   K�
   V�   a�   l�   w�   ��   ��   ��   ��   ��    ��   ��   ��    ��   ��   ��   ��   �   �                            ������    ��   ��   ��"�   �                               "�   @                       ������    ��   �   ������   '�   2�   =�����H�   S�	   ^�
   i�   t�   �   ��   ��   ��   ��                    "�                          �����    �   &�   1�   <�   G�   R�   ]�   h�   s�����~�
   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �   �                        "�                          ������    ��   ��   ��   ��   ��   ��   ��   ��   ��������
   ��   �   �   �   %�   0�   ;�   F�   Q�                    "�D   �                       ������    ��   ��   ��   ��   ��   �   ������   #�	   .�
   9�   D�   O�   Z�   e�   p�   {�   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ������
�   �    �    +�!   6�"   A�#   L�$   W�%   b�&   m�'   x�(   ��)   ��*   ��+   ��,   ��-   ��.   ��/   ��0   ��1   ��2   ��3   ��4   �5   �6   �7   (�8   3�9   >�:   I�����T�<   _�=   j�>   u�?   ��@   ��A   ��B   ��                                                            "�    \                       ������    ��   ��   ��������   ��   ��   ��   ��   ��	   ��
   	�   �   �   *�   5�����@�   K�   V�   a�   l�   w�   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��                                "�   �                       ����p�    {�   ��   ��   ��   ��   ��   ��   ��   ��������
   ��   ��   ��   
�   �    �   +�   6�   A�   L�   W�   b�   m�                        "�G   �                       ������    ��   ��   ��    	�   �   �   '�   2�   =�   H�   S�   ^�   i�   t�   �   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �   �   �   $�   /�   :�    E�!   P�"   [�#   f�$   q�%   |�&   ��'   ��(   ��)   ��   ��+   ��,   ��-   ��   ��/   ��0   ��1    �   �   �4   !�5   ,�   7�7   B�8   M�9   X�   c�;   n�<   y�=   ��>   ��   ��   ��A   ��   ��C   ��D   ��E   ��                                                            ������"�   "                               �    �"    �����"�   T"                              �"`���        D    ����    ,   ��        �    �"    ����@�"�   �"                              #`���        ,D    ����    ,   ��    ����    ����    ����    `#    ����    ����    ����    <    ����    l���    ����    �C    ����    ����    ����f0f    ����    ����    ����    +g    ����    ����    ����    �v    ����    ����    ����    D{    ����    ����    ����    �~        W~        ����    ����    ����    0�    ����    ����    ����    ҇    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    &�    ����    ����    ����    ��    ����    ����    ����    ա    ����    ����    ����    F�    ����    ����    ����    ��    ����    ����    ����    `�    ����    ����    ����    [�    ����    ����    ����    *�    ����    ����    ����4�:�    ����    ����    ��������        Θ    &       $&��        �H    ����       ��        ����    ����    ����    ��    ����        ����    ����    ����    X�    Y�f�        ����    ����    ��������    ����    ����    ����5�;�    ����    ����    ����#�.�    ����    ����    ��������    ����    ����    ����o�|�    ����    ����    ������    ����    ����    ��������    @           N�����    ����                  �'"�   �'   �'                       ����    ����    ����    P�����    ��        ����    ����    ����    ������    �        ����    ����    ����	��    ����    ����    ��������    ����    ����    ����    �!    ����    ����    ����    �#    ����    ����    ����    .%    ����    ����    ����    u'    ����    ����    ����    �(    ����    ����    �����*�*    ����    ����    ����    �1    ����    ����    ����    �=        e<        ����    |��    ����    I        zF        ����    ����    ����    �V    ����    ����    ����    �]    ����    ����    ����    ]a    ����    ����    ����    Ld    ����    ����    ����    ��        ��        ����    ����    ����    c�    ����    ����    ����    !�    ����    d���    ����?�E�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    r�    ����    ����    ����    �    ����    ����    ����    q�    ����    ����    ����    8�    ����    ����    ����    ��    ����    ����    ����    O�    ����    ����    ����    ¾    ����    ����    ����    ��    ����    ����    ����    >�    ����    ����    ����    x�    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    !�    ����    ����    ����    ��    ������"�   �,                           ����    ����    ����        ����    ����    ����    �    ����    ����    ����    �����    -        ����    ����    ����    r����    �        ����    ����    ����    p        \        =            ����    x���    ����    �b    ����    x���    ����    Sd    ������"�   (.                           ����    ����    ����f    ����    ����    ����Yksk    ����    ����    ����    e�    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    8�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����g �     �����"�   �/                           ����    ����    ����    �
    ����@�"�   (0                           ����    ����    ����    A:    ����    ����    ����    R<    ����    ����    ����    ?    ����    ����    ����    �J    ����    ����    ����    �S    ����    ����    ����    V    ����    ����    ����    �X    ����    ����    ����    W\    ����p�"�   X1                           ������"�   �1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       6ڀL    9          �8 �8  9 3� 9   vrmlexporter.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ||�Y    .?AVLODObject@@     �Y    .?AVObjectData@@        �Y    .?AVNodeData@@      �Y    .?AVBaseData@@      �  �Y    .?AVbad_alloc@std@@         �Y    .?AVexception@std@@         �Y    .?AVlength_error@std@@          �Y    .?AVlogic_error@std@@       |�Y    .?AVNavigationInfoObject@@          |�Y    .?AVStartDialog@@       �Y    .?AVGeModalDialog@@         �Y    .?AVGeDialog@@      �Y    .?AVVRMLSaverData@@         �Y    .?AVSceneSaverData@@        �Y    .?AVConfirmTextureCopyDLG@@         +  8  d  ||||||8   |||||||||�  �Y    .?AVDisjointNgonMesh@@          �Y    .?AVGeSortAndSearch@@       �Y    .?AVNeighbor@@      |||   ||?  �  |�Y    .?AVGeUserArea@@        �Y    .?AVSubDialog@@     �Y    .?AViCustomGui@@        ||||�Y    .?AVTexturePreview@@        |||   v   �   �Y    .?AVResourceDataTypeClass@@         |D   g   �   |||l   |����||||�Y    .?AVout_of_range@std@@          �Y    .?AVinvalid_argument@std@@          N�@���Du�  s�      |�Y    .?AVtype_info@@         |�Y    .?AVbad_cast@std@@      �Y    .?AVbad_typeid@std@@        �Y    .?AV__non_rtti_object@std@@         PZ              �?pow     acos            sqrt            cos             sin             fmod         4rF�߈F���F�߈F�݈݈�݈F�F�߈F�                       �|    �|                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����   ��������                       |�Y    .?AVbad_exception@std@@                     ��������    ��������������������        |�                                                                                                                                                                                                                                                                                                                                                 ����         ������������                                         	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                             ۋ               ��       ���ܧ׹�fq�@      ��@�6C����?      �?exp          !�����a�                             ���5�h!����?      �?                         �   P	   
   h   0   �   �   �   \   ,   �   �   �   X   �    �!   x"   �x   �y   �z   ��   ��   �                                        �����
                                                                      ?           x   
       �D�D                       
      p?  �?   _       
          �?      �C      �;      �?      �?      ���d�j�o�u�z�������������ɏΏ�����>�C�]�b�����������&�:�R�f���������ʑޑ��
�*�/�I�N�n�������ΒӒ���&�>�R�r�w�������ʓ�                                                                          H!                                                                                                                                                                                                                                                                                                                                        abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     �P�  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                                                                                                                                                                                                                                                            ������C                                                                                              �V            �V            �V            �V            �V                              �\        �� ��� \�V   �V�P                                                |l �                              �      ���������              �        �p     ����    PST                                                             PDT                                                             0XpX                                ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l                      ����        ����                                                                                                                                                                                                                                                                        �&     �+   �+   �+   �+   ��   ��!   ��   �+   �+   �+   |�   t�   �+   �+    �+   �+   �+   l�   �+   d�   \�   T�   L�   D�"   @�#   <�$   8�%   0�&    �                                                       �D        � 0             ����           ����    t�p�l�h�d�`�\�T�L�@�4�(� ������ �����������ح̭ĭ�� �������������t�p�l�`�H�<�	                                              \.   �\DwDwDwDwDwDwDwDwDw�\               .                         ���5      @   �  �   ����                         ��������             �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (�         �� T�                     �� �� �� ʔ Ҕ � � � 4� L� X� j� ~� �� �� ̕ �� �� �  � .� F� `� ~� �� �� ��  Җ � �� 
� � (� >� T� `� r� �� �� �� �� �� ȗ ؗ �  � �  � ,� B� R� h� v� �� �� �� Ę ֘ � �� � � 6� P� j� x� �� �� �� �� ʙ �� �� � � "� .� <� L� V� b� n� �� �� �� �� ؚ � � � (� 8� D� T� j� z� �� �� �� �� қ � �� �  � 2�                                                                                                                                 �� �� �� ʔ Ҕ � � � 4� L� X� j� ~� �� �� ̕ �� �� �  � .� F� `� ~� �� �� ��  Җ � �� 
� � (� >� T� `� r� �� �� �� �� �� ȗ ؗ �  � �  � ,� B� R� h� v� �� �� �� Ę ֘ � �� � � 6� P� j� x� �� �� �� �� ʙ �� �� � � "� .� <� L� V� b� n� �� �� �� �� ؚ � � � (� 8� D� T� j� z� �� �� �� �� қ � �� �  � 2�                                                                                                                                 ` CopyFileA KERNEL32.dll  �InterlockedIncrement  �InterlockedDecrement  !Sleep �InterlockedExchange �InitializeCriticalSection � DeleteCriticalSection � EnterCriticalSection  �LeaveCriticalSection  �RtlUnwind ZRaiseException  -TerminateProcess  �GetCurrentProcess >UnhandledExceptionFilter  SetUnhandledExceptionFilter �IsDebuggerPresent �GetModuleFileNameW  OGetSystemTimeAsFileTime �GetLastError  C CloseHandle FileTimeToSystemTime  FileTimeToLocalFileTime �GetFileInformationByHandle  >PeekNamedPipe �GetFileType l CreateDirectoryA  FindFirstFileA  .FindNextFileA �GetCurrentThreadId  oGetCommandLineA �HeapValidate  �IsBadReadPtr  � DebugBreak  zWideCharToMultiByte MultiByteToWideChar �lstrlenA   GetProcAddress  �LoadLibraryA  4TlsGetValue �GetModuleHandleW  2TlsAlloc  5TlsSetValue 3TlsFree �SetLastError  �GetCurrentThread  �GetModuleHandleA  FatalAppExitA ;GetStdHandle  �WriteFile :OutputDebugStringA  �WriteConsoleW ;OutputDebugStringW  ExitProcess �SetConsoleCtrlHandler �LoadLibraryW  �GetModuleFileNameA  �SetStdHandle  �SetHandleCount  9GetStartupInfoA x CreateFileA  CreateFileW JFreeEnvironmentStringsA �GetEnvironmentStrings KFreeEnvironmentStringsW �GetEnvironmentStringsW  �HeapDestroy �HeapCreate  �HeapFree  WVirtualFree TQueryPerformanceCounter fGetTickCount  �GetCurrentProcessId AFlushFileBuffers  �GetConsoleCP  �GetConsoleMode  �HeapAlloc �HeapSize  �HeapReAlloc TVirtualAlloc  RGetACP  GetOEMCP  [GetCPInfo �IsValidCodePage #GetProcessHeap  \VirtualQuery  LFreeLibrary �InitializeCriticalSectionAndSpinCount kGetTimeZoneInformation  �GetLocaleInfoW  �GetLocaleInfoA  �SetFilePointer  �SetEndOfFile  hReadFile  �WriteConsoleA �GetConsoleOutputCP  �LCMapStringA  �LCMapStringW  =GetStringTypeA  @GetStringTypeW  hGetTimeFormatA  �GetDateFormatA  �IsValidLocale � EnumSystemLocalesA  mGetUserDefaultLCID  R CompareStringA  U CompareStringW  �SetEnvironmentVariableA                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        <   L5�5�5Z6�6�6�6�7�7;8�89f9�97;h;t;�;�;v=�=�=>>�>�>  8   �0�0M1�1�1�1�1s2�2�23/3�9�9�9�;<�<�<d=�=�?�?     $   �5�5�7q9�9�9�9�9�9�9�9 :�<{? 0 @   O0�0O1�1�1�3�3808<8H8T8`8?9�9�:�:�:�<�</=`=l=�=k>�>�>   @ d   1-1~1�1�1�1�1�1�23�3�3�4�4n5�5�5�5,686D6P6\6�78{9�9l:�:�:;#;i;�;�;*<d<p<_=f=�=>6>�>�?   P 4   �0�0T1�1�2�2�3�3V44�6�6�7�7<8A8�<�>?�?�?   ` h   00�0 1�1242@24(4446<6H6�8�8�8�8�8�8�8�9�9�9�9�9�9�9V::�:;$;�;�;�;�;<<"<�<==(=D=I=N=   p <   �0�0�1�2�2�2�2�34/4V4�5(6�6�6*7�7�7v8�8�8F9o9:;i<   �    /0f6�6T7&8P8E9Y9�=   � �   (0�273P3\35/5f5P6l6v6�6�6�6�67797C7d7z7�7�7�78$8,8084888<8@8D8H8L8P8T8f:�:�:�:�:�:�:!;+;O;Y;z;�;�;�;�;�;�;�;�;�; <<<<<�>F?m?�?   � `   0�0�0�0$1o1�12*2@2V2l2(5>5�5�5�67�7�7�8�889D9P9h9l9p9t9x98<�<=#=i=�=�=*>d>p>�>?�?�? � <   0�1�2�2�2�2@667]7�7�7�78 999�: ;;X;d;p;o=�=�>�>   � 0   [0�1�56 6,686V:}:�:�:�;�;�;�;�>�>�>�>   � 8   �1�1�122�5�5 666$606<6�92:B;H;�; <,<�<�<�=   � P   0I0�0�0�0 11:1�122�2�2P3 4f5�5�6�9�:4<l<x<�<�<�<�<�<�<�<�<�<�<r?�?�? � \   90�1�1�1�5�57<7H7T7`7l7x7�7�7�7�7�7�7�7�7�7�7�788 86;_;�;�;<===�=�=�>�>(?4?�?�?   P   80=0N0
1D1P1\1�12;2@2Q2�2 33v3�3�5�5f9�9�9�9:?;p;|;�;6<_<-=`=l=b>??    4   V00�3�3�304<4�45�8�89�9�9�;�;�;�<�<�=�=        i2�2�2�4�4�6�6v>�>�? 0 L   00&2O2�23&4O4�4�4f6�6778H8T83:X:d:�;�;==,=8=T=Y=^=|=�=�=�=�= @ H   �1�1�1�1�1�1�1�34$4f5�566_6�6�6v7�7�7�7�:�:�:�; <�<=4=@=�>?   P L   �0�0�0�4�4�5�5�5�5�5�5�5�6�6�6�6�6�6�6f7�7�7(848�8�8 99(9-929�=�=   ` @   �01.2�2�23?366_67/788�8�8�8�8�9�9�9�9v<�<F=p=�=�=f? p <   �0�1�1�1�1�3�3�3V77�7�7�7�7�7-929C9O9k9p9u9�<�>�>   � @   X1h3�3�3g8�8�8�8�89[:�:�:�:�:�;�;�;�<�<�<'=@=L=?�?�?�? � H   �0�0.1V2}2�36-6�7�7'9@9L9�94:�:�:�:;�;-<f<�<�<�<�<f>�>�> ??   � ,   1%1�1�1�1�7�709�:�<�<�<==�>�>H?^? � X   0E0j0"1T1y1�1�1b23y3�3P4�4*5�5�5�56�8�879M9�9::a;�;�;�;�;�;X?e?q?~?�?�?�?   � X   �0�1�1212M2v2�3$4�4�45�5�5^6�6�6�7�7�78�8�8�89=9j9\:�:;,;B;X;�>�>�>?�?�?�? � D   1H1T1`1l1x1�1R8�8�8P9u9�9�9�9�9�:;0;`;l;x;�;|<T>�>�>�>?�? � 4   0+01n1�1�144f4�4f6�6�67-7C7�9�9�9�9=?=? � D   0-0Z0�01$1�3�34*4�6�67c7�7�7�9:�:�:�:n<=�=�>�>?$?:?P?  	 (   �4�4%6>6T6j6�6�6�6�6_=�=	>">8>�? 	 H   0(040@0L0X0d0p0|0�0�0�0�09F9l9x96:]:�:�:;><W<m<�<?'?=?S?i?    	 ,   �2f5�586�6�6�69*9@9V9i<�>�>�>?�?   0	 @   �0Y3�3�3�334?4M4�4�46(6>6*7@7V7l7
: :6:L:�< =�=>??   @	 <   L0b0^1t1�2�3�324H425_5�5�56 6,686D6P6=�=$>Y>�>�>   P	 d   �0m2r2{2�2�3Z4�455�56-6B6�677 7�78-8B8�8Y9�9�9�9?:M:b:�:b;�;(<4<@<�<="=�=">�>9?h?t?�? `	 T   f0�0202<2H2T2�3�3�3�3�3_4�4&5�56�6747�718�8(9Z9�9_:�:K;�;?<�<?=�=?>n>�>�? p	 X   0�0E12�2x34;4�4�4�4�4`5�56g6�6�6�6/7�7{89�9:�: ;G;l;x;�;b<�<b=�=b>�>b?�?   �	 <   b0�0G2�2G3�3�425�58�8�8�8$909�9R:�:�;2<�<r=u>?�?   �	 H   ?0�0B12�2�2k3�3K4�4+5�56{6�6[7�7r8�8�9::;�;(<�<�<f=�=Z>f?�? �	 @   0�0�0P1�12E2�23Z3 414�4�4�5�5
6�6�6\7�7:�: ;�;<�<�< �	 h   =1G1Q1[1e1o1y1�1�1�1�1�1�1�1�1�1�2�2 3O4�4/5�56�6�6h7�7878h8t8�8b9�9K:�:2;�;;<�<=�=>�>;?�?   �	 H   0�01�12�23�3�3o4�4b5�5a6�6a7k8�8�8�;<<=<=H=I>l>x>{?�?�?   �	 8   �0�0�0�172�2�3 4,4:5`5l5z6�6�6�7�7�7:>`>l>{?�?�? �	 @   �0�0�064�45o5�5V6�67�7"8�8;9�9":�:;�;<�<�=�=:>l>x>�> �	 P   0{0�0k1�1O2�2?3�3�5�5�5�5"6�67�78�89�9:�:+;9<\<h<t<�=�=�=�=M>�>*?�?  
    O04�;`<  
 <   �415`5l5�5n6�6�627�7/8�8B9�9O:�:R;�;?<�<1=�=!>�>!?�? 0
 D   "0�01�233�3�45{5�5[6�6;7�778�8+9�9:�;Q<�<k=�=[>�>Y?�?   @
 <   K01�12�23{3�3�4�4�56�6�6�78�8;;@;Q;�;�;�;<<< P
 8   '0�3�3�34404b5g556:6r7�7�7�7�7�7�78888r<R= `
 <   1�1�4�4k5�5K6�6N7�7�8�89E9�9�:�:�:�:M;�;R<�<|=�=v> p
 @   �0�0�0�0q1�3~4�4v5x7�7�78�89x9]:�:h;<�<*=�=>�>?�?   �
 @   0�01�12{2�2_3�3�465�5�667�7k8�8[9�9Y:5<�<�<�<�< ==   �
 P   0�0/1�1224u4�4�4�4R5�5�677�7�:�<�<�<�<3>B>Q>b>q>�>�>�>s?�?�?�?�?�?�? �
 h   82�2�3T4�4d5�5F6�67�7�7o8�8�8�8�89�9�9:(:4:�:�:�: ;,;�;�;<@<L<X<�<�<&=3=�=�=>,>>2?`?l?�?   �
 \   30�0�0?1\1�1�2(3�3C4�4N5�5J6�6*7�78�8�89;9h9t9�9::�:�:m;�;F<�<M=�=>�>??�?�?�?   �
 `   00�0�0f1�1/2�2�2f3�3F4�4:5�56,6b6�6�6�6j7�7]8�8*9�9:o:�:�:�:�:O;�;-<�<8=�=>�>�>m?�? �
 `   J0�0&1�12v2�2!3D3P3\3h3�3444@4L4X4�45$505<5H5�5S6C7/8�8;9�9;:�:;�;<v<�<?=�=>�>?�? �
 `   0 1$101�12�2
3}34�45v56�6!7�7?8o8u8�8�8�899�9O:�:�: ;_;�;<<<�<(=4=�=>H>T>�>M?�? �
 T   @0�0&1�12}2�2O3�3J4�45�56�6�6m7�7�8V9�9/:�:/;T;`;�;<�<�<k=�=>->�>�>K?�?   h   ;0�071�12-2�2�2�2�2?3�314M4�4�4�4�4Q5m5�5�5�56�6k7�7_8�8_9�9O:p:�:�:�:?;�;?<�<B=�=/>�>??�?    P   �0�0o1�1r2�2r3�3[4�4?5�5?6�6?7�7?8�8?9�9�:�:�:;D;P;\;�;a<�<�<=�=�=�=     8   �5�5	6�6�6�6�7p8�8p9�9r:�:r;�;_<�<8=�=.>�>U?�?   0 d   H0�0;1�12�2�2o3�3]4�415M5�5�5�5�5Z6�6:7�78�8�8f9�9?:Q:�:�:�:�:O;a;�;�;�;�;j<�<�<�=�>6?�?   @ H   ;0�01�12�23�34�45�56�67�78�89�9":�:;�;R<�<`=�=`>�>_?�? P L   b0�0d1�1_2�2_3�3_4�4_5�5o6�6r7�7_8�8`9�9[:�:K;�;+<�<"=�=:>�>�>,?�?�? ` @   00�3�3�3�4 5�56�6 7�748�8�849d9p9|9�9�:�:{;�<�=L>�>�? p 8   ;0�0�1+2Q3H4x4�45�5�586h6t6<�<�<�<C?I?�?�?�?   � \   �0`1�1�1�1P2�2I4�4�4 5�5Q6�6�6�6�7F8l8x8�8$909�9�9�9�:�:�:1;�;�;�;!<u<�<�<j=�=�=�=   � 8   A6T6M8|8�8J:�:�:�:;;[<�<�<=�=�=>$>�>Z?|?�?�? � �   J0l0�0�041�1282D2�23(343�3�34$4�4�455�5P6r6�6�6@7b7�7�708R8x8�8 9B9h9t9:0:X:d:�: ;H;T;�;<8<D<�< =(=4=�=�=>$>�>�>??�?   � \   `0�0�0�0N1p1�1�1>2`2�2�2/3	404<4H4T4�4�5�5�56�6#7�738�8N9�9n:�:~;!<�<,=L=�=r>?�?   � @   G0�0a1�1�12(2�2n34�4J5�56�607�7P8�8v9:�:T;�;�<�>�?   � T   �2�3�3�3�3�3 4444�4$6(6,6064686<6@6D6h8H9`9�9z:�:�:^;�;><�<.=�=M>�>Q?�?   � L   a0�0�12�23~3�4$505<5H5T5`5l5!6�6&7�78�89�9(:�:m;�;^<�<f=
>�>�?   � ,   ?011�1J2�26D7#9b:�:�:�:�<�=�>f?�?         o0�0Q1�1�12�2�6/7�768�8  P   �1�1�1�1�1�1�1�1�4!5O7t7�7+8P8\8�8'9X9d9M:t:�:];�;�;n<�<�<�=>>?<?H?�?      k0�0�001H5p5|5�:�:�: 0 \   40474>4E4L4t4�4�475Y5`5g5n5u5|5�5�5�5�6�6�6�6 7�7�788:�:�:k;�;_<�<_=�=D>�>$?�?   @ L   0{0�0;1�1+2�23�34�45�56�67�7K8�8/9�9:|:�:P;�;0<�<=�= >{>�>r? P H   t0�0_1�1J2�2�2�2�2�2s3�3�3�56�677�78�8a9�9�9�9�9_:�:K;�;�>   ` P   
0�0�01<1H1�1K2�2+3�34�45�5R6�6o7�7o8�8o9�9r:�:X;�;H<�<8=�=(>�>?�?   p 4   0�0�0�1�1�1*2�23�3;4`4l4�4�67�7�7�=�=t>y> � `   �1�1�1�1�1�1�12222)232=2G2Q2[2e2o2y2�2�2�2�2�2�2�2�2�2343@3 4b8u88�8�8�8�8�8�8�8   � 4   �8�8�89 9)9?;D;M;�;�;�; =%=.={=�=�=�=�=�=   � ,   p1�1�1�1�2�2�5�5�5�5�5�5�5�::=`=l=   �    0�0�0�0 �    ~4�4�4'6L6X6�67_9   � P   �2`3d3h3l3p3�4X5�5K6�6/7�7/8�89�9':�:;�;<�<=�=>$>0>?D?P?\?h?t?�?   � H   X0�0g1223�34�45�56�67�7+8�8;9�97:�:/;�;<�<=�=+>�>�>�?   � `   0�01�3Z4�4�428X8d8V9^9�9�9�9�92:7:@:�:�:�:�:�:�:�:5;\;`;d;h;l;p;�<�=�=�=L?R?z?�?�?�?     �   00E0w0}0�0�0#1k1�1�1�1/2_2�2�2�3�3�3�3�3�3�34L4]455'585X5�5�5�5�5J6n6�677(7H7�7�7J8t8�8�89+9K9k9�;�;x<>>? ?%?  x   �2�2�2�23333333#3)3-33373=3A3G3K3Q3U3�3�3�3�5�5�5�6�6.7�7^8�8>:�:�:*;N;�;�;<Z<�<�<=7=�=�>�>�>�>�>n?�?�?   �   h0m00�0�0�0�0�01(1R1W1\1�12'202~2�2�2�2�233&3N3�4 50555:5?5�5�5�5�5+676V6p6|6�6�6�6�6�6�6�6
767R7^7n7z7�7�7	888F8K8P8U8|8�;�;�;�;�;B<K<u<z<<�<�<�<�<�<�=�=�=�=�=>>A>F>K>o>x>�>�>�>2?r? 0 �   *070G0T0?1�1�1�2�2�2�2�233L3U33�3�3�4�4�455�5`6�6"7�7�7�7	88�8�899/9w9�9�9:8:=:O:�:�:�:�:�:�:";:;C;x;};�;�;�;�;�<===P=u=�=�=�=>%>Z>_>d>�>�>�>!?&?+?Q?i?r?�?�?�?�? @ �   00C0M0.181�1�1�1�1V2h2�2�2W3i3N7X7�7�7�78	8868?8l8q8v8�8�8�8�8�899J9Q9�9�9 :<:@:D:;>;J;z;;�;�;�;�;�;�;<+<[<`<e<�<�<�<�<v={=�=�=�=�=�>�> P p   �0D2H2L2P2T2�4�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::::: :$:(:,:0:4:8:<:@:D:�=
>#>�>�>�>�>2?r?�?�?�?   ` �   010<0N0�0�0Y1g1y1�1�1�1�1q2v2�2�2�2�23
33b3�3�3�3�4�4�4�45,5�5�5�56�6�6�6y7�7
8@8�8�8\9~9�9�9�9*:_:x::�:�:�:�:�:�:;;;;;;; ;$;n;t;x;|;�;�;�;<<<< <A<k<�<�<�<�<�<�<�<�<�<
=====�>�>�>�>�>�>�>(?-?2?   p �   �0�0�0�0�0p1�1�12!2+282l2}2�2p3z3�3 4(4-4?4e4n4�4�4�4�4�4�455\5h5�5�5�5�5666f7x7�7�7�7�7�7�7�7�7�7�7�7�7&8/8b8~8�8�89.9X9a9k9�9�9:!:=:[:�:�:�:�:==/=x=�=�=�=�=�=>->\>3?   � �   �0�0�0�0�011 161B1K1P1Y1e1n1�1�1�1�1�12e2j2�2�233'3/383@3F3L3T3Z3`3h3y3�3�3�3�34�5�5666E6h7m778�8�8�8�8�8�8�8�8�8�8�8999V9[9�9�9:/:4:U:u:�:�:;;S;a;�;�;�;<	<<<&<.<;<D<J<S<X<^<f<l<�<�< ==P=Z=f=�=�=�=�=�=�=�=�=�=>�?�?   � �   00011/1U1a1�1�1�1�2�2�2(30393I3U3k3w3�3�3�3�3444B4N4�4�4�4�4$5*5b5h5�5�5�56"6[6g6�6�6�6�6�6�6%7/7;7V7s7}7�7�7�7�7h9m99�9�9�9�9�9�9:: :,:B:N:W:}:�:�:�:�;�;�;�;<<�<=#=F=�=�=�=�=B>G>L>l>q>�>�>�>�>�>�>?j?v??�?�? � �   0_0�0�0�0!1r1�1�1�1 22(3-3?3S3�3�3�3�3�3�3�34!4'444�4�4�455>5C5H5X5u5�6�6�6�6�677/7	8'939V9h9m99�9�9�9�9�9:K:�:;;;F;#</<\<a<f<�<�<�<�<�<�<=.=3=8=�=9?J?b?s?   � �   h0m00�0�0�011j1z1�1�1212C2[2�2�263;394+5\5a5f5�5b6r6w6�6�6$7)7.7]7y7�7�7�9�9�9�9�9:+:X:]:b:�:I<f<�<�<�<�<="='=e=q=�=�=�=]>�?�?�?�?�? � �   11@1]1�1�1�12�2�2�2�2�2�3�3�3�3.4�4�4�4�4B5�5�5�5/6O6t6�6�6�6�7�7�7�7\8g8�8�8 9%9�9�9�9�9�9�9�9�9::::&:F:O:X:e:s:�:L;S;�;�;�;,<`<e<�<==9=?=E=i=o=u=�=�=�=�=�=>>   �     p1}1�5�5J6�9�9�9�<�<�<   � 4   H0M0_0X3]3o3�4�4�4�<�<�<(=-=?=�=�=�=h>m>>   �   00m0�0�2�2�2�2�2�2�2�23l3�3�3�3�3�3�344(4�4�4�4�4�4�4�455O5y5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�56666 6&6,61666<6A6G6P6W6^6s6�6�6�6�6�6�6�6�6�6�6�67+727^7888'818:8A8G8x8}8�8�8�8�8�8�8�8 9>9�9*:2:O:s:y:�:�:H;M;_;><{<�<�<�<�=�=�=�=�=>>>1>;>B>w>�>�>�>�>�>�>�?�?�?�?     �   <0B0H0N0T0Z0a0h0o0v0}0�0�0�0�0�0�0�0�0�0�0�0�0�0�01111/161�1�1�1�1�1I2O2]2g2	6T6`6�6�6�6�6�6�6�6�6^8j8�8�8�8�8�8999X9d9�9�9�9w:|:�:�:{;b=n=�=�=�=�=�=>>>V>b>�>�>�>  H   �6D7P7}7�7�7�7�7�7�7�739?9l9q9v9�9�9�9�9�9)<x<�<�<�<�<�<�<==#=   �   �0�0�0�0�021<1�1�182=2O2u2z24393>3H4M4_4�4�4�4�4�5�5�5�5�5l6�6�6 788/88:=:O:;a;j;�;�;�;�;�;&</<Y<^<c<�<�<=A=J=t=y=~=�=�=�>?,?6?N?e?�?�?�?�? 0   0-0:0G0T0�0�0�0�0�01M1�1;2b2i2�2�2�2�233H3M3R3�3�3�3�3�3�3�34�4�4�4�4�455$5.5>5H5W5�5�5�5�5�56�6�6�6�6�67!7<7I7N7T7a7f7l7�7�7�7(8-82878j8v8�8�8�8�8�8�8�89999C9H9M9R9�9�9�9�9#:(:-:2:]:b:g:�:�:�:;;;;9;B;t;�;<�<�<�<==%=7=A=_=d=i=�=�=   @ �   00601	11"1'1O1U1p1}1�1�1�1�1�1222R2W2\2a2�2�2�2�2�2�2�2�2$353:3?3D3m3r3w3|3�3444M4R4W4\4�4�4�4�4�4�45!5&5+5N5W5�5 6�6�6�6 777S7Z7i7�7�7�788J8Q8[8m8w8�8�8�899�;<�<�<�<�<=�=�=�=�=�=E>u>�>~?�?�?�? P   
0b1l1�1�1�1�1�1222#2+2C23W3�3�3�3�3�3�344/494G4L4S4]4a4k4z4~4�4�4�4�4505=5I5Y5u5�56K6P6]6b6p6�6�6y77�7�7�7�8�8�9�9�9�9�9�9�9:0:5:::R:�:�:�:�:�:;';3;`;e;j;�;�;�;�;�;<</<�<�<�<�<�<�<=	=,=3=V=^=�=�=�=	>>>;>A>�>�>�>??G?L?Q?x?|?�?�?�?�?�? ` �   �0�0�0�01�1�1�1?2F2M2j2�2�23)3V3[3`3�344�4�4�4�4�4�4�5�566�6�6�6�6�6777-727<7J7O7Y7m7s7{7�7�7�7�7�7�7#8.8Q8\8}8a9m9�9�9�9�9�9:	::�>�>�>�>�>??J?S?}?�?�?   p �   00A0j0s0�0�0�0�0�0Z2�2�2�2�2�2�2�2�231383<3@3D3H3L3P3T3�3�3�3�3�34!4<4C4H4L4P4q4�4�4�4�4�4�4�4�4�4�4:5@5D5H5L5w6�6�6�6�6�6�6,757@7{7�7�7�7�7�7�7�7888`8�8�89Y9e9}9�9�9�9A:�:�:/;7;�;�;�;�;�;�;?<l<�<==�=�=�=	>y>�>�>?�?�?�?�? � `   0M1z1�1�1D5�5�5686U6i6t6�6�708�8L9�:�;�;�;�;�;�;�<�<�<.=�=�=�=�>�>7?@?j?o?t?�?�?�?�?   � �   !0&0+0T0]0�0�0�0�0�0�0�0�0?1H1r1w1|1�1�1�1�1�1C2L2v2{2�2�2�2�2�2 32393�3�3�3�34G4S4�4�4�4�4�4;8c89"9L9Q9V9�9�9�9�9�9N:S:X:v:{:�:�:�:�: � �   r1z1�1�1�12%2H2c23,3@3P3\3e3�3�3�3	4�4�4�4�4�4�4�4D6L6q6y6$8�8�8�8 9939>9W9`9|9�9�9�9�9�9�9�9�9�9/:4:9:@:m:r:w:|:�:�:�:�:�:�:�:�:�;�;<x<�<=I=N=S=�=F>Y?x?}?�?�? � �   
0"0�0�01/1W1]1f1{1�1�23363D3R3h3�34%414X4d4p4�4'5J5V5�5�5�5�5�5�566$6G6�6�6�617@7�7�78*8F8{8�8x9}9�9�9D:O:�:�:�:�:;2;q;�;�;�;�<�<�<�<�<�<�<�=�=G>�>�>m?t?   � �   �0�01+191L1�2�2�24442474<4]4b4g4�5�5�5:6C6m6r6w6 77�7�7�788E8J8O8�8�8�8�8�8�89/94999�9�9�:�:�:�;�;<<#<T<[<�<�<= =%=> >M>R>W>�>a?�?�?�?   � t   0<0^0h0�0�0�0�0�0u1�1�133q4-5�56�6�6$8L8x8�8�8�8 9S9b9�9�9�9�9�9�9 :::�:�:�:�:�:�:�:�:�:�:x?}?�?�?�?�? � �   00�0�0X1]1o1�1�1�1�1�122J2O2T2�2�2�2�2�2=3_3�4�4�4p5|5�5�5�5�5�5r6~6�6�6�6�7�7�7�7�78�8I9l9�9�9�9�9�9:H:j:t:�:;&;G;�<�<>�>�?�?   � �   +070�1�1	222a2�2�2�2�2363p3�3�3�3�3�3�34444 4$4(4,404449$9*9Y9$:,:A:�:�:�:�:;O;�;�;3<p<�<�<=_=�=�=>c>�>�>?W?b?�?�?   �   00k0v0�0�0#1o1z1�12c2�23l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3T4X4\4`4d4h4l4p4t4x4|4�4n7�7)959E9Q9n9t9�9�9�9�9~:I;U;e;q;�;�;�;�;<<�<�<�<Z=n=�=�=�=�=6>Z>i>~>�>�>�>�>�>q??�?�?�?�?�?�?�?  �   0e0m0�085A5P5\5g5q5�5�5�56@6c6q6z6�6�67$7�7�7�7�7�78X8]8c8t8z8�8�8�8�8�89&959<9L9U9\9b9i9o9�9�9�9�9:#:0:8:G:\:h:t:�:�:�:<<<�=�=�?�?   l   k1w1�12\3�3�3444�4�4�4�4:5F5v5{5�5�5�5�566�6�67�7�7�7�7�7q8x8�9�9�:�:�;j<�<w=�=�=�=�=�>?L?�? 0 L   555555 5$5(5,5054585<5T5X5\5`5d5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 @ �   <01&1V1[1`1�1�1:2L2�2�2�2�2�23)3Y3^3c3�4�4 66<6A6F6�6�6$7)7.7|78(8X8]8b8-949E:Q:�:�:�:|;�;�;�;�;)=5=e=j=o=`>l>�>�>�>j?q? P �   �0�01�1�1�1�1�2�2�2�2�2�3�3444�4�4 5%5*566J6O6T67*7Z7_7d7�799J9O9T9:*:Z:_:d:�:Q;<<O<T<Y<#=/=_=d=i=>>@>E>J>6?B?r?w?|?   ` �   90E0u0z00$1�1�12#2(2^2j2�203q3�4�4.5358566>6C6H6&727b7g7l768B8r8w8|8i9u9�9�9�9y:�:�:�:�:�;�;�;�;�;�<�<�<�<�<�=�=>
>>�>�>???�?�? p �   +00050�01;1@1E1�6�6�6�6�6w7�8�8�8�8�8\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::::: :$:`:d:h:l:p:t:x:|:   � (   4;q;�;�<�<�<�<�<�<h>�>�>�>�>8?`? � 0   e6�7�78�8�8�89a:|:�:q;{;�;??H?�?�?�?�? � �    0
0G0�0�0�1�1�1�1�12 2%233A3F3K3q3z3�3�3�3�3�3
444�4�4�7�7�7�7�788=8O8�8�8�8�8�8�899�9�9�9:):2:\:a:f:�:�:�:�:�:�:;7;A;z;�;X<]<o<�<�<�<===B=Z=c=�=�=�=�=$>->?T?]?�?�?�?�?�?�?   � x   4090>0d0�0�0�01o1�1�1�1�1�1�2�2E3y3�3�3�3�34b4�4�4�5�5(6D7N7x7�8�8�8�89t9~9�9�9=A=^=�=�=�=>X>]>o>�><?�?�?   � �   00$0e0l0�0�0�011>1C1H1o1x1�1�1�1�1^2w2�2�2333)3d3m3v3�305n5~5�5�5�5�5�5�5�5v6�6�6�6�6�6�677797I7U7�7�7�7�7�7 8&8T8Y8^8�8�8�8�8�8(:-:?:e:n:�:�:�:�:;t;{;�;�;�;�;�;<�<�<�<�<===*=<=B=�=�=�=
>U>??�?�?�?�? � �   >0�0�0�0�01(2-2?2f2�2�2�23
33�3�3�3�344"4�4�4�4�4�4�45"5+5A5Q5k5t5�5�5�5�5�5!6-6Z6_6d6y66A7M7z77�7�7�7�7�7�7�78{8�8�8�8�8�8�8�8 9%9*9B9�9�9�9�9�9�9�9�9�9�9:":+:H?U?^?x?�?�?�?�?�?�?�?�?�?�?�? � l   000(0/050>0D0O0Y0h0q0z0�0�0�0�0*232�2�2�2�2,383Y3�377 7�8�8�8�8�8�8�8�8�8�8�89959S9Z9�9�9�:   � �   �3�3�3�3�3�3�3�344"4.4?4K4T4`4h4t4{4�4�4�4�4�4�4�4�4-5=5g5X;];o;�;�;�;�;�;<<�<�<�<=r=�=�=�=�=�=�=)>X>�>�>�>�>�>�>�>�>�>�?�?   T   #030=0b0l0�091�1�142�2�23L4t5{5�5�5�5�5�5�6�67%7�;�;�;�;<g=�=O>[>�?�?�?�?  �   050[0�0�0121N1j1�1�1�1	2!2�2�2�2�2�2�3^4�4�4�4�4�4�455 5$5x5}5�5�5�5�5�5�586=6O6�6�678?8�8�8�:�:�:�:�;(<-<?<�<�<�<�<�<=�=�=�=>>>F?O?U?]?c?o?t?�?�?�?�?�?�?�?�?   T   �0191b1�1�1�1�4�5&6+606�7W8�829H9^9x;�;�;<<<<�<�<�<�<g=}=�=�=�>�?�?�?�? 0 x   �0�0�0�0Y1^1c1�2�2�2:3?3D3�3�3�3�3*4/444�4�4�4}5�5�5�5�5Q6Z6�6�6�6�6�6�6�6�6�:�:;;7=C=�=�=#>,>9>C>K>P>W>�>x?? @ X   00�011&1-1@1^1c1�1�1�1�152J2u2�2�2�3=4I4�4�4�4�5�5�5�5�5'78�8�9�:�;w<g=W>G? P T   '0(4�4�5i7�89-92979\9e9�9�9�9�9�9:::::C:m:r:w:)<�<�<�<�>�>�>???%?V?   ` �   �1�1�1K2{2�3�3�34<4�4�4�4�4�4�4555&5/555�5�5�5�5�5�5�5�5-626�6�6�6�6�6�6�6�6 777�7<8I8r8|8�8�8�8�8�8�8�8999t9�9�9�9�9:3:�:�:�:�:�:A;F<T<x<�<�<�<�<==1=V=_=h=s=|=�=�=�=�=�=�=�=�=�=�=�=D>c>p>�>�>�>?
??2?E? p    J0Y0b0�0�0�0�01;1C1I1m11�1�1 222-252[2b2h2q2�2�2�2�2�2�2393D3[3f3�3�3�34D4R4a4j4�4�5�5�566*636X6`6y6�6�6�6
777"797D7S7y7�7�7�78P8T8X8\8`8d8h8�8�8�8�8�8�8�8�8�8�8�8�8�8`9d9h9l9p9t9x9�;�;<<<!<><G<i<u<�<�<�<�<�<�<�<H=Y=l=w=�=�=�= >>7>>>D>S>a>i>�>�>�>�> ?4?E?`?s?�?�?   � �   +0o0�0�0�0�0�0�12%2.2�2�2�2�2�2�2�23'303[3n3w3�3�3�3�34E4M4X4`4h4�56 6-6<6E6^6l66�6�6�6�6�6�6�6<7J7k7t7z7�7�7�7�7�7�7�7�7E8�8�8�8�8�8�8i9�9�9�9�9�9�9::*:7:?:D:W:d:s:|:�:�:�:
;-;:;|;�;�;�;�<�<�<�<�<�<�<�<=	=4=e>�>�>�>�>�? � <   G0P0�0�0�0�0�0�0�0�0�0�0�0 111�5�5�9-:�;1<W<d<�>�? � 0   q0+1T2f35�5�627�7�7�=�=�=�=�=�=	>>_?   � �   00#0)0C0J0�0�0�0�0�0�01111(11171E1R1[1d1�1�1�1�1�1�1�12292�3�3�3�3�3�3�3$4m6{6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6P7T7X7\7`7�7�7�7�7�7�7�7�7�7�:�:�:�:�:;�;�;�;�;�;�;<:<�<�<�<�<.=5=�=�=�=�=�= >>v>�>�>�>"?+?<?W?n?w?   � 4  A0[0b0�0�0�0�0�0+141:1T1[1`1h1�1�1�1�1$2(2,20242|2�2�2�2�2�3�3�3�3�3�3�3�34O4W4g4p4�4�4X5j5�5�5�5�5�5�566(6?6�6�6�6�6-7X7�7�7�7�788!838E8W8i8{8�8�8�8�8�8�8�8	99-9?9Q9c9v99�9�9�9 :::&:�:�:�:�:�:�: ;�;�;�;�;<<@<D<H<L<P<T<X<\<`<d<�<�<�<�<�<�<�<�<�<�<�<�<=== =D=H=�>??'?.?4?=?B?W?f?u?�?�?�? � �   000 0$0(0,000A1R1q1v1�1�1�1�1�1�1�1�12D2H2L2P2T2X2\2`2d2h2�2333>3L3T3`3l3{3�3	4#4�4�4�4�4�5)8:8H8U8�9�9�9>:F:y:�:�:�:�:�:�:�:;;f;s;{;�;�;�;�<�<�<�<n>w>}>�>�>�> ?	?�?�? � l   R0w0�0�0�0O1x195P5^5g5x5�5�5�5�5�5+6�6I7s7j8';@;I;N;�;<)<F<W<�<�<�<�<�<�<	== =E>r>�>�>�>�?�?�?�?   � 0   0&0F0f0�0�0�0�01&1T1b1�1�1$2466<Y<�=        �4t7M89[:�>  T   F1�1�2�34�4�4�6�7g8�8�8�8�8 9	99#9/9;9^9e9�9U<a<m=�=>>/>V>�>)?2?\?a?f?     �   *0R0B1�1G3O3�3�34"4'4h4p4�4�45$5)5�5�586@6}6�6�6�6�6a8j8�8�8�8�8�8&9/9Y9^9c9�9�9:1:::d:i:n:�:�:;?;H;r;w;|;�;�;!=*=T=Y=^=�=�=�=�=�=[?�?   0 �   "0.0[0`0e0�0�0�0�0�01F1N1�1�1�1�1�1 2'2Y3e3�3�3�3�3�3+40454w4�4�4+5�5�5�5�5+60656r6z6�7]8+949^9c9h9�9�9�9�9�9::N:W:�:�:�:�:�:�:;;�;�;
<<<Q>]>�>�>�>�>�>�>�>�>5?=?�?�?�?�?�?   @ �   00;0@0E0;1G1t1y1~1	3F3O3y3~3�3�495m5�5+7�9�9:::V:^:�:�:�:;	;i;q;�;�;4<@<m<r<w<�=�=>>>c>k>�>�>�>�>�>\?d?�?�?�?�?�?�? P �   q0x0�0�0�0111K1S1�2�2�2�2�213=3j3o3t3k5�526>6k6p6u6�6�6�6�6�67X7_7�7�7�7�7�738;8i9u9�9�9�9::;:@:E:�:�:�:A;�;�;<<G<L<Q<�<�<+>�>[?d?�?�?�?�?�?�?�?�?   ` �   50=0�0�0�0�0�0�011161;122G2L2Q2�4�4�4�4�4	55B5G5L5�5�5�5�5666V6b6�6�6�6�7�7�7�7�7�:�:�:�:�;<=<F<p<u<z<�<�<�<�<===,=6=h=q=�=�=�=�=�=�=�= >�>5?A?q?v?{?�?�?�?�? p x   0�0�01�1�1�2�2�3�3�4�56�6�6777�7o8�8�8\>`>d>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???????? ?$? � D   A5M5z55�5�5�5�5�5�5�7�788$8�8�8 9R9�9�9�: ;;;;;;;; � �   0O0�6�6�6�6�6�697B7l7q7v7�7�7�7888-8�8�8�8�8�899B9G9L9�9�9�9�9�9�9:�:�:�:�:�:�:;$;>;K;S;�;�;�;H<M<_<�<�<�<�<�<�<===@=J=S=X=]=�=�=�=�=�=�=�=�=�=�=�=>	>4>@>s>>�>�>�>�>�>??6?;?@?Z?�?�?�?   � �   111(3-3?3�3�3�344)474B4J4R4Z4d4l4t4�4�4�4�4�4�4�4�4�4�4�455525:5B5J5R5^566 6.6C6Q6k6y6�6�6�6�6�6G8V8/9>9�9�9�9�9�9�9:":':,:P:V:]:g:m:v:~:�:�:�:�:�:�;�;�;�;�;<<E<J<O<f>o>   � �   �0�01 1%1a1j1�1�1�1�2�2[4;5G5N5x5�5�5�5�5	6&6^6j6p6�6�6�6�6�6�6�6�6�6�6�6777%73797D7N7`7�7�7�7�78*939]9b9g9�9�9::Q:Z:�:�:�:�:;�;�;�;<<:<?<D<�<�<G>�>�>�>�>�>??(?3?d?�?   � �   0(0"1.1�1�1�1"2E2N2�2�2�2�2�2�2333R3�3�3�4�455H5f5�5�5�56;6D6y6~6�6�6�6�6777L7U7�7�7�7�7�78�9�9�:�:;B;x<}<�<�<�<�<2=7=<=b=z=�=�=�=�=�=�='>,>1>j>�>�>�?   � �   0$0\0a0f0�0�0�0�0�0�01%1]1b1g1�1�1�122262s22�2�2�2�2Y3}3�3�3�3�34*4X4�4�4�4!5E5k5�5�5�5�5g6�6�6�67H7h7�7f8p8z8�8�8�9�97:[:�:�:;';`;�;�;�;�;4<T<r<]=g=q=�=>4>S> � �   �2�2�213T3]3�3�3�3�3�3�344"4[4�4�4�5�5�5�5*6H6�6�6�677?7D7I7�7�7�7�7�7�788(8R8W8\8�8�8�8�9�9s:�:�:�:�:
;);J;d;�;�;�;�;�; ==9=>=C=[=a=�=�=�=�=�=>W>�>?�? � 8   �0/1�5167777�9�9�9:%:0:S:^:�:>>b?w?�?�?     |   00070L0�01H1�1�1�6�6�7�7�7�7�7�8�8�89999*909P9�9�9�9�9�9::":)<4<F<]<�<�<�<=/=4=9=�=�=>>>�>�>??5?:???  8   77M7�7�7�7�78#8(8�8�8�8�8�8�=�=|>�>�>!?&?+?�?�?   `   00Z0f0�0�0�0�0�01#1(1�12N2Z2�2�2�2�2P3\3�3�3�3@4G4U5\5�6�6n798�8F9R9�9�9�9g:�:;S;   0 �   �0�0'1,111�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12222 2$2(2,2024282<2@2D2H2h9m99�9�9�9�9�9�:�:;
;;�;�;<�<�<�<�<�<�<�<==&=0=K=R=[=r=y=�=�=�=,>8>p>u>z>�?�?   @ `   �0S1�2�2�2�2�23B3K3�3�45T5�5*6R6�607Z7�7�9�9�9�9:::$:�:�:/;�;�;�<�<�<=�=�=�=�=�=   P ,   �9):s:s;~;�;�;�;�;�;%<�=>1>�>�>?   ` X   �1"2>2S2_2�2�4�45%5D5c5�5�5f6|6�6�6�6R7z9�9�:;;B;P;^;=,=�=�=>,>~>�>M?�?�?�? p �   000�1�122b2g2l2�4B5G5L5�5�5�5,61666�6�6�6�6�67]7b7g7�7�7�7#8(8-8�8�8�8; ;M;R;W;�;�;�;�;�;<<E<J<O<�<�<===�=�=�>�>�>??   � �   �0�0�0�0�01	1m1y1�1�1�12!2N2S2X2�2�2�2�2 34�4�4�4�4&525_5d5i5�5�5666�6�6�6�6�6<7H7u7z77�7�78$8)8�8�8�8�8�8]9i9�9�9�9::E:J:O:�:�:�:�:�:];i;�;�;�;<<E<J<O<e=q=�=�=�=)>5>b>g>l>?'?L?P?T?X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�? � P   �6�6V8]8|8�8�9�99:E:;;<$<$=0=�=�=�=�=�=�=�=�=�=�=�=4>8><>@>D>H>L>P>   � 8   ~0�0�0�34�4�4T5Y5^5c5�5�5�7�7<8�8�8�:�=�=,>~>   � <   E0K0�0�0�1	2#2K2X2n2}2�2C3|3�3�56�6�7�7�7}8�8�8�8   � $   �2�:�;a<m<�<�<�<6=a>h>�?�?   � @   �0�0�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 666H6L6P6I9S9w9Y: � `   Y0�0!2&2+202�2�2�2�2�2�2�2�23!3&3+3�9%:1:a:f:k:�:�:�:�:�:�;�;<'<W<\<a<�<8=?=N>U>�?�?   � p   m061�1i2u2�2�2�2�34?4v4::J:O:T:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;4;8;<;@;D;H;L;P;T;X;\;`;d;h;l;     \   �4�5�5�5�5 6E6Q6�6�6�6�78*969f9k9p9::N:S:X:�:|;�;�<�<�<�<�<�=�=
>>>{?�?�?�?�?    �   �0�0�0�0�0�1�10373�3�3�344�4�4555i6u6�6�6�6{7�7�7�7�768h9t9�9�9�9z:�:�:�:�:7;�;�<�<�<�<�<�=�=�=�=�=�>�>�>�>�>�?�?     �   000�0�0111�1s22�2�2�2�2�2�3�34�5�5�5�5�5�6�6�6�6�6�7�7�788�8�8999::A:F:K:;#;S;X;];0<<<l<q<v<B=N=~=�=�=i>u>�>�>�>{?�?�?�?�?   0 �   �0�0�0�0�0�1�1�1�1�1&727b7g7l7829>9n9s9x9�9�9�9�9�9�9�9�9�9 :::::(:,:0:4:8:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: @ (   (:-:?:e:n:�:�:�:i;�;�;4<@<==�? P �   �0)1�2�2�2�2�2333E3N3x3}3�3I4R4h4�45#5�5�5�5k6w6�6�6�677;7@7E7�7�7�7�8�8�8[9g9�9�9�9�9�9::":�:�:�:h;m;;�;�;�;�;�;�<=2=`=�=�=>�>�>�>�>	?�?�?   ` �   E0K0P0u0{0�0�0�0�0�0�0�0�0�0�01i1�1�12�2�233M3g4p4�4�4�4�4�4555�677;7@7E7n7w7�7�7�7a8j8�8�8�8�8�8999G9P9z99�9
;(;4;a;f;k;�;�;�;�;�; <<9<><C<�<�>�>??]?f?�?�?�?�? p @   00050:0�5�576M6�6�6�6�67#7(7�7�7�7�7�7<<�<�<!>->�>�> � X   �0�0�0�0�0'101Z1_1d1�1�1�1�1�1�3�3�3�315):4:>:E:O:Y:e:p:�:�:�;�;`<�<�<�=$>J>�>�> � �   11G1L1Q1�1�1�1�1�1�12-22272�3*434]4b4g4�4�4551575?5M5S5f5�5�5�5�5�5�5�5666#656A6�6�67]7m7�7�78!8&8�8:q:�:�:Q;z;;�;G<P<z<<�<4?:?@?F?L?R?X?^?d?j?p?v?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? � �    000000$0*00060<0B0H0N0T0Z0`0f0l0r0x0~0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�011111 1&1,12181>1D1J1P1V1\1b1h1n1t1z1�1�1�1�1�1�1�1�1�1;2}2�2�2l3�45[5�56@6�67r7�7�7-8|8�8L9�9�9:E:�:�:�:;M;};�;�;"<�=�>�>�? � L   �0�2�3�4#6�6�67~7�7*8�8�89k9�9�93:�: ;�;�;-<~<�<=w=�=->|>�>1?u?�? � @   0l0#1u1�1�1T2�2�2M3�3�3)4�4�45Y5�5�56]6�6v81:�:�;-=q> � (   �14�59�9*:Z:�:�:�:�:�:*;Z;�;�; �    �<�<A=v=�=   �    �=>6>    `   1222 5$5(5,505@8D8L9P?T?X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?     014181<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222|2�2�2::::: :�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<\<`<d<h<l<D=H=L=P=T=X=\=`=d=h= ?$?(?,?0?4?8?<?@?D?H?L?P?T?X?\?`?d?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? 0    00000 0$0(0,000 P �   d4h4p4t4|4�4�4�4�4t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6064686<6@6D6H6L6P6T6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7�7�7�7�7�7�7�7�7�7�7�8�8�89 9$9�9�9�9�9�9�9�9 : :$:(:0:4:8:@:D:H:�:�:�:   `    �?�?�?�?�?   � (   l9p9t9x9|9�9�=�=�=�=�=P?d?h?l?   �    (0,0 P 0   l6p6t6�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< p �   �7�7�7�7 88888888 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8d8h8l8p8t8x8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99999999 9$9(9,9094989<9@9D9H9L9P9T9X9\9`9d9h9l9\=`=d=l=p=t=|=�=�=�=�=�=�=�=�=�=�=�= � �   �2�2�2�2�2�2�2�2�2�2 3333 3(30383@3H3P3X3`3h3p3x3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 4444 4(40484@4H4P4X4`4h4p4x4�4�4�4�4�4�4�4 5(50585@5H5P5X5`5h5p5x5�5�5�5�5�5�5�5�5�5�5�5 � �  33$3,3034383@3X3d3|3�3�3�3�3�3�3�3�3�3�34 4(4<4@4T4X4l4p4�4�4�4�4�4�4�4�4�455 5(5,50585P5\5t5�5�5�5�5�5�5�5�5�5�5�5�5�56(6,6@6H6L6P6X6p6|6�6�6�6�6�6�6�6�677$7,7074787@7X7d7|7�7�7�7�7�7�7�7�7�7�7�7�7 880848H8P8T8\8t8�8�8�8�8�8�8�8�8�899$9<9@9T9X9l9p9�9�9�9�9�9�9�9�9�9�9 :: :8:<:P:X:\:`:h:�:�:�:�:�:�:�:�:�:�:;;; ;8;P;T;h;p;t;x;�;�;�;�;�;�;�;�;�;�;<<(<0<8<P<h<l<�<�<�<�<�<�<�<�<�<�<�< == =8=<=P=X=\=`=h=�=�=�=�=�=�=�=�= � �  004080<0@0D0H0L0P0T0X0\0`0d0h0l0p0t0x0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�6�6�6�6�6 7747@7d7p7�7�7�7�7�7�7 888808P8X8`8h8p8x8�8�8�8�8�8�8�8�8�8�8�8�8�8�89949<9H9p9x9�9�9�9�9�9�9�9:,:L:T:\:d:l:t:�:�:�:�:�:�:�:;;;@;H;T;X;d;x;�;�;�;�;�;�;<<<@<H<P<\<�<�<�<�<�<�<=(=0=P=X=d=�=�=�=�=�=�= >>0>4>8>D>X>d>x>�>�>�>�>�>�>? ?D?P?t?�?�?�?�?�?   `  0(0@0H0T0�0�0�0�0�0�0�0�0�0�0�0�0�0 1111 1(10181@1H1P1X1`1h1p1x1�1�1�1�1�1�1�1�1�1�122$202\2|2�2�2�2�2�2�2�2�2�2�2�23333$3,343<3D3L3T3\3d3l3�3�3�3�3�3�3�3�3�3�3�3�3 4444 4(40484@4H4P4X4`4h4p4x4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 50585@5L5x5�5�5�5�5�5�5�5�5�5�5�5�5�5 6666 6(60686@6H6P6X6|6�6�6�6�6�6�6�6�6�6�6�6�6�67777$7,7H7T7x7�7�7�7�7�7�7�7 8(848\8|8�8�8�8�8�8�8�8�8�8�8 990989@9H9T9|9�9�9�9�9�9�9�9$:,:4:@:h:p:x:�:�:�:�:�:;;; ;(;0;8;@;H;\;h;�;�;�;�;�;�;�;<<8<@<L<t<|<�<�<�<�<�<�<�<�<== =D=L=X=�=�=�=�=�=�=�=�=�=>>(>L>X>`>�>�>�>�>�>�>�>�>�>?? ?L?l?t?|?�?�?�?�?�?�?�?    �  0040@0h0�0�0�0�0�0�0�0�0�0�0,1<1H1P1t1�1�1�1�1�1�12,242<2D2L2\2h2�2�2�2�2�2�2�2�2�23,3P3\3d3�3�3�3�3�3�3�3404T4`4h4�4�4�4�4�4�4�4�450585@5H5P5X5`5h5p5x5�5�5�5�5�5�5�5�5�5�5�5 6666 6(60686@6H6P6X6`6h6p6x6�6�6�6�6�6�6�6�6�6 7777 7(70787@7H7P7X7`7h7p7x7�7�7�7�7�7�7�7�7�7�7�7�7$8D8L8T8\8d8l8t8|8�8�8�8�8�8�8�8�8�8�8�8999$9,949<9D9L9T9\9d9l9t9|9�9�9�9�9�9�9�9�9�9�9::: :(:0:8:@:H:P:X:`:h:p:x:�:�:�:�:�:�:�:�:�:�: ;;;; ;(;0;8;@;H;P;X;`;h;p;x;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<< <(<0<8<@<H<P<X<`<h<p<x<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<@=`=h=p=x=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>> >(>0>8>@>H>P>X>�>�>�>�>�>�>�>�>�>�>�>�>�>????$?,?4?<?D?L?T?\?�?�?�?�?�?�?�?�?�?�?�?�?�?   �   0000 0(00080@0H0P0X0`0h0p0x0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 1111 1(10181@1H1P1X1`1h1p1x1�1�1�1�1�1�1�1�1�1�1�12 2D2L2X2d2�2�2�2�2�2�2�2�2�2 3333(3H3h3�3�3�3�3�34(444X4x4�4�4�4�4585X5x5�5�5�5�5�5�56666(6<6`6h6l6�6�6�6�6�6�6�6�6 77 7<7@7\7`7|7�7�7�7�7�7 8808<8\8`8|8�8�8�8�8 9 9<9@9`9�9�9�9�9�9 : :@:`:l:�:�:�:�:�:;0;P;p;�;�;�;�;<0<P<p<�<�<�<�<�< =@=`=l=�=�=�=�=�= > >,>8>l>p>�>�>�>�>�>?0?P?p?�?�?�?�?�?�?   0 (    0,080p0�0�0�0�0101P1\1h1�1�1   @ �   000$0D0`0�0�0�0�011D1H1h1�1�1�1�1(2,2024282<2D2H2L2P2T2X2\2`2d2l2�2�2�2�2�2�2�2�2�2343T3X3\3`3d3�3�3�3�3�3�3�3�3�3�3�3�3 44,4l4p4�4�4�4�45p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�8�8<9@9D9H9L9P9T9X9\9`9l9p9�<
====t=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>$>�>�>.?2?6?:?>?B?F?J?N?R?V?Z?^?b?f?j?n?r?v?z?~?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? P �   00
000000"0&0*0x0�4�67 707@7P7t7�7�7�7�7�7�7�7�7�8�8�:�:�:�:�:�:�:�:�:�:�:;;;;$;,;4;<;D;L;T;\;d;l;t;|;�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ====                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        